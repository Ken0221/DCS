`define CYCLE_TIME 5.5
`define NUMBER_OF_PAT 10
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
cpsqx1Xq4Wy0IxW1uiZ/rCjV7fDi8QndlTFueNS8JlvQHC6/HiFuuSa01NbMcYkD
64YHhvXr8pImbOItZWPZz3jPsdDyR2Ug6Trz7LOdvvqa3BKNp+sNfT6zyNXd1vXN
RRs+lRkpCOp6wf6RhN5NeWVMYsrF4pMGx0pp/eouHOynUK99tEnL6rRh+JZSnPzH
c+6EJsGriRFeGducTkgrCxRN2P6pNPqLWpZ6xHh9iThRvHEwOPMbxxOXT7Ssgm0I
YF9K/VAOvehS/g34L/IHjvuqCqaleR+hyAvM27Wrd+O+I4ih6nOV78ZSRN3oBQsz
1cenDQA5dyHroUdrAYMXHg==
//pragma protect end_key_block
//pragma protect digest_block
/9szycdIRlzhtP1qG03XVpNVSD8=
//pragma protect end_digest_block
//pragma protect data_block
iticwMI8trXa+VnRf2bthZdRFctkg4HcJF/kxNT/VQWf6npGL60r4mOiIUqnfVxL
dsoSQdFq8F6jCynbp7XNmznR04pJIe6Md7NRiOCtCgjyBmxVjVA0hna/2mJar3rK
gJkrwqLbZT7HIhYGB0KISbQXX3B2WgHUW3BQt5V5KC8b5TIuGTq1Ao3GOooq+1tb
WfAsAvX/8ER33Flz/a2XiaDauSXyvUQIpaLuS96PR1JagFOkzNTsXyEm5+w0ykAL
SAmGNugKKghzNZzy5NJEjFlMGb2Da+DegoIJSDJv5j5h3uuWWJFW/ZMRwjsWqTY0
BU3GRI+3t4YF+V24jlQo91gEIr4CYJqoDRaArXVOzj2lneNo7JEWhfEhtDetyl+4
wxaog1uAkOI8V0xw2Iv5gGlwqtp7zB+4JuFkVNoZcn+go2fX797GMIoRJ8lEWcdj
F1r3VXuavCOSzSccxw+DdXkBZv5nfE7z8A+CY8aUnkA+Jm82Ni+eDAHpYn0LUCzI
baRsDzUp89RH1IO/CRcJCcATZ8SZfz6buYZgmBExfP9ofXNq6D31KPb3VR6Sr3sC
daaje+C0DdM/gksvcKuwIU1BDENiGvITVfDULNPlFCc88VdIIMSamuJEvOKliuLa
ArVbbX3F9ilrR1bAGlKe7SrSx0Kmf/PJR4ll0LVW5i1yo9gY0q6VPWH08H9BOuEw
w26mtCY7RCsrFwv5mwOtxhUj38Qrpvt+WA9vLOaGOgGDVrA2CAlGbMDtOzbDYeem
StSFcsXktmjMfgZxb/SNbbV48iZVxsCOtyKgHOSU1c4k7/lKz2mO2DKlmSlOIVo/
ACIxpmIexPsmKMJu6vgNytEDdLfruBPuv/PfsylprRr7227/R0cBkAYTqLKS/2ZN
sM/4TWVJH6lPKY7n46reod1DWbf5CEe+IgOjTE+N+6GYK7rIaXkwQENov35iYiHA
rbsUVrkFjzqSYI/wJMTJcBF8Dkjn75gVPYywaFMMSbevOB2GdRJGSKuG1VEDN2jn
/w/YDoSUFIEloZBlrMn+hgDNohF1QtsezV3cPHyiTCPIQZWbtTVJvU7mDYXTU5Ka
TWlGhsbso81F65iYTwXRs+vHjGFgwqY7vzdsT85QhH1t1eUlFTA2w99HxxE8/0nc
q1qzbfUI72KPAmWZ4DLmLL21I2wJmARFbnxBOptjd9Y3EXkuHUzdNKRzCeKEm0HP
YsmyrYJd2AduHLOqN//erbnqpK2C4MkGgxAftazHFcvXG9p7LshnzR93JcnXPguL
oFNzhbC32I58dlZQy2nA9RBcESu57rbEGHT10PkbPhvryYWen+KYl/2qtW4xHRid
jLW8t6Tc+NVk7kYNYVHFxx9Oh/EuuY2K85w2YrkIygd81YEyPttQJigtXBX0rq+j
2QF7gdLmKM7gc4u845cv8m52Vxa8uqSQuJeXPnqk3mN7RJoI5p/zbmIIiNehhipZ
Pe27fWskJ+70emqlQLd5OcQx/Lzyaqw54zZpekPtYLrJ504/1zXfExKceCWj4tvP
SCIZ1yw5wiXgOwzv6ZBbpE++1XEDPwKn2PyA8Bs6AJru5lSPADjMOsB2Tk8pv7QR
pzB+r+l13Aocse9x+GXOAerIWe0O2BrMkkZMau9sW5AG/jKjA7+ZfDqnkvgwhPsh
AvsM6GDCNQIJaI0EAG/CU4+VM4W6dKSLFK8wag/M/SjPAaSgSYit4QEQ26z5f3m9
u/6Irt2BsaATTGRKa1/MkaBkRQOeqDcKw/woo5pq61wervxewYiR/0PRYWBs9CrY
3LB82N499kFu2BL9g0LRdEKa8ncw2erIYL6cl6/1+RQXvUHsCWKRHHTukQcQ/sKF
Z/Spg3GGC4F160afzQXC6Sys40oqMbCa++LjpnC/axgES8S6JTVwom7s8a+1L/UC
t4VPBeuFCHlrwU4oSboovai6Zz27QB8ppyN4py2ZxYrI15duWx73Jw2NYFdGqIW6
tWfGGzsE6LuGOsDji8LGphrCXtZ4g/HoFd0Lq2ikK+RV6f13mxDzbIt4OkP+2KCp
VgCbXIfusPshacWo+AI3dQhoEUbQc8TPfI+WgzfSJiWJli2fS0oiXyMOan6XAGE5
5pqNOc+qHgn4LsOZtoxtrEAv9PWZg7gjACfMHKKY8elIS9iw/D1fCU8bpb35g3m+
EN+KGwaHZPqAVghaH2D3omPpOIVhEygWZaLDjJ6GmuburmhQPVzgNah+bQe1ug9L
mgyeQyvg/RAJ9Hg8FxkflwtTueaduTq0rvu64j+GIf9mcHnZ67U6wrmv0rrhfd9h
fj+XfQPBhQSJywtE2jzf6uTfSyjzo2Qc2CP40hyLEjgJDxwr6iqBR09Z1+bt3maU
ZcjkvPhFzx3ghLxBjg7BaOzYz0bfO1gJepzpON13Y+lH3i9evrek6fUs8DuFCr+G
unGFK/2dlMCvWCYqPTSf3yPxL/IRcAc/Ffe4+JPoPKlGwjA5uIKCtWiU8JA1QIbp
z94sn7jeHbsOQVMaWgN7OzEDYmpmbYQHL0NZFUltBw6YIVyTI5rLiwBPVImCVemB
+enVFzMB4tGwcV1okt24WqI8RRKpDSkgWPA9PA9nglkjZdKL2scn3jG2EZpdmkN6
Ai/e377W+OJusbRMzklqFC75o8GeODCUwmGZQG/mNbkuY/nrF5paoVhuTodpcJmk
/S9KaTCjYSU+GtQPnWWugNvN9i7RSMj1MT4QfC8hX0rPzq0pjUvQvE7ypl0XImmK
Ua+M6STUzPoXwajcnKxrzcy9xc+GlSRdNZXMJxcl8fcbQOcos2ZY4na7zVkxU7jt
9A3Kza64roideNRz2LJ91bx27oLym5sqSMzEcSlekySgYUNE/HFKBywSCNiG9DmQ
zm/IaKsa7jnAHjZp3Mse6qIuleBvkGYzqBmhHo51O3gGF/RGqBL1u5Au6vcDKBNL
RyLRV6ZsmGHQ9vtjgYCDmWasHtwWgbS/fFzgH/k86HXRjSTAKHresWN5o6BqtvaE
CqtluNroF2sGLJxSkQrM47joM7e9AgYqDOvxKQd1MyUqspRq19/SxOxPzFsHv7v3
c4byh83qzZ4VxDku5WsTWwO3IfOKur6275mJqUzyxjC0s+1epM+OhECT5rScTHcr
pLQ7eY3+flaRQ/m2u8v2b73XOG6kky2zmXHkEbpkVX1vTHVVeE9mAxbAvrcNZU9o
LrTZ+Cmzj9RFNqWlWqlyMv226e3GqNlp4OZHPJf0AU/KY8J/+Fibot+DuwiYNUl9
+yCtHk0pOejcBhT1jDeR5K44uxZeZteGQBc/EMQuufxcpr1eqeL19pJBBmXXuZmZ
BV4PgfJkkXNC87Dflp649hYpk2M+nLOF/nCuwRGf4LyGv5owrb0sM4ChNQU4t8Zl
CaiaSRQ3WrpIzQ4wfAKOL3g4XUyluFmK9foghvj0dworyGltoV7iWJCdcJ4qByE0
Z29lUk//A6Kz16O6Y9Cxjy43fCuIJSkT53STbcxdmZufA+8DBTXB0/fBLILAOO3v
gOtiuOMzKPWzShYPQwlkHjdm8T08eS66JE+b/D7hGSXZP/dHauh0l2lYhHHHmSC0
8qM1rxmVNv3yNBHxinQod/tCNeGWm681ptSkNesfhTStDBej5Jja1EATLilBmile
lR1uXSffIgw3fx3yHi0uULsv0peNHDQBHm+qiEG8flS/R0kDf/KmtGTnC7ZInnPN
5fYDMZhGG9XNhqfJvAxhhmC7407VlJqpJN3P0pTwijRBvJgUk00Usn0WIPuA7YHp
nfVQNGCfUlu9i26p4+L2jbi4LD5BLLKlzxpbhMwoCHrrjGRW9RaS6ab5f3aY8Soq
eAmb79xrW1pGk9xLSq4ykPGVxVCKq2QXYAdICSl7qq1KvedoDrs35AT1BCN9x7zG
acJr5j4VnkJQpRhDF61k7AnPgqWWs5Gqn2f9eLSqU3AT79S0y1eEGj+65G2zxW40
TBdAD1dyDdCc3M6YH+EG+WPXQmhWUPv64NST3L3FxJ7jBiD+1RvVUv+mH8GSBXvo
ZlXk+h5FCkSAfYEyo5v1VJd8d5Zv0fpLbFivdw9p5snGutNBweTMtqQUm8PZWouB
AE6YHi29rq8IwoV3NrKOB+DBxF3FpO3dgU4IgWmXNC3bTDw66vciay+PA9wdqPza
2hgrnSyoe2ym6PpNvZOZ5TgGa04Jpeaw0DjevtXgp327H7tNTJJjUMC7CFzOfrA9
BAat2Shyql1B5Rr56UaZvK+xH9PX2Fh93HCCrnU1T+IJj/M4YtYsVV2YY1YMkUkv
YOFcrTE/7Ljy8I2KYtCyqNUOeLMT9JxNMBYEXo07GelrtDOSKjZtYLM8e8PLmUbL
TJL8XRpkQ0EYJpKvc9XGUQTD76hl+/XysX0HGVVb0228aqDrrOZ2ClMF1DGwKRc+
pTS5DvJE5TCXjSyR+MKByxgFaw7OY+R3+yNVHWYGzrdWR3IiHNOLJtFfR51RUtiP
aoSHHjaob6ZO+tLAk437qMVUccXfOrick80YlP8VY8G0CcDOZC3xKw2pOkJLbrX5
bQHU5Fl6MbwtO4OM4C3Ni4u9+uYqMEc6q9MthXGEEEd0KFLvHR8ETwCPr+Nnve2h
YFlOtIsX9aANvzhkaBdnOSUlmJUxgw1OIXhAHqhshCmLcWb1hyYRSbMFcORVayqv
kALBVsMkObIo4okfWXKHKSy7SOw9QJSVXTkT0KQ5Zm8h2l2F6rzITezXmA6Kfpde
SLN7qD7qsk1OppXG6HZBCkt9cPFnEYJyGqWr8xIw4M4ePC4/QgMH0k01mvTqP1d/
o4qQYeiKUk/g3nl/95QmzHU08CGUNo3BDsbunlRCkgjxGyTV08BSQ9OEJn9N9awd
psUoieNU44eFG9eCU6QpoiosEv90zdI6tw+5f+6RiBTYMYoGDe/ZiBXnvxOdc8sf
PPDK/yYfcDcV9SSZLzvxrcN+w9Xjg49dWTf4GCYFwl0pEB/U9MZPtRj0eYkdvqQz
gMRfzYdPUh72oeOSX7b2/vwmI91gu7OZG5eI/rQUFXAhRzNXAQZB6X1Qr9RKKitW
GWNsgLxd2n3Ft1ZiGlPL2iInJYVKMJ2V6utByVPZBQXj80hZsx6YZZ2SXe0sRwgb
cLq8T+8Kv05pxlbqfzUIJZNcCJvEUtpAlAQt5FncMQYqYPmcjGlNdBYLVeO4Zor4
6p9NOnXiu6kEv+R9Ac+bLqoocMXJWI9gV3DXTDB1oRiXXOa6LogWmelJxr+YJtZv
lSqXwkMD/scNPLcngD6lhvGhLALFAtRnWaifmt9K5WYJRiOIq5TjSKBmfWnrY5Ol
JVCS8nnnY54sTku6ELbuA7W+ML9ThXNGVoHzI+GC9e8sTIUvbHuOUKkf/U+uxb6C
JDduIcYV016266CXOdD8hNjryrPIEXShSoReoHWLoTWjEu8Q3MaGfI/3cwKU2VaT
za5BUTIJQkjhJJZ+WTSzjsSlPGC7Wi1UQdUQ8yy6rcQn6ji4ux/mIuyL9PQNeMnx
6mxbcC4Kj06OLh0l+6xJ2Bs16EHsCX3H0Sb305vvLMlENr7HKx7wWdL6LkvVt+/m
s8/+tr7+ZaclTE8MI2nUMBwiaGjqCjC1IG3nXWvHwFzK8OI1R+KIYFkCgzwfs7Mo
TfuG48zkZ90uDc8vJIawweEAxGuRyb6BQRioIihgnuuvLEpJksjGae8gjuS2PAss
7xLBVWcS4mp2j+N7GyDk8KXwBmNCtQMJtTXc1+g7aife3nOk7dVxSluSA3XEyaSc
6FTuXnhoSKHHYZZzBPoOHlgKVSSRBsvY4bkb2oAtPRZmBo99aY6Qwe4whlb2kbuH
usowSDChhn8ShhSoDlwFICJeqluKT6YUjK1SExXaenDZKiuG0tmVHZ9kCxhRr6Q2
YYpJSo53ulPTq9lItMN2Zo3mbh2rSGzkTz7nDqGrH2kq+o3NuZvdvh5qP1u5eEKh
P4WhTBIDoYQYJ1uYdGymCqNaEQVsIFWXS9rai9goHnqYOtWatzgV3r5KvLX4H+aD
z4H/nWniaY8jR6Xa6WGP/VDdsNaBG+f3fYmSJsfCnwTnsBN7BjEmgUHhXgFhoj5G
KGt3NMDQ/fbMEgwsdEwLU1qu3yfU/LGd4E6Xe+NyocetxV+o1EopGbHquBHU5AoS
UN1MZbeRMeR694uADoQi8Qji6rXEYmW8tM2d26t7t1ORcGjVVSketoO7xsPAVanx
klupa/rysnHh+Ku1PFZDL00AH2gHaRJPrgOnamj+GE+ExMMzyy6mq8FAjmEu4cPr
wcwyCxtTpOSt4QykLBihJH/gHedq4Z3019l0iex+4uJch6BvlJdeKhfJTcFgS0bC
GGcgYf47lfWtUsz4JK7A0IIIvK1oYu10GhU6h56RrWwoKb1RmS68FtD1ocmxawov
U0WZUnVBLQGlwVG50MF/hWPKaxnZmEHliYy49rgfSyhLRJ6vKIln2fBGq6iiLSjQ
wMOMRrNfs34RQVlZyhd+pNzpvhv6ZmrBPclG0wyVyi1R9e2TZbw4b+rVP1dHrN8N
GCLDS5AEj1dNaDW1KsDxRvkXnPcVK3oyrGg6tOhiP+XhyaT3tPDd2hDH2TlLzH1o
6iEElxDLYtLhtKhEQhU4pGdPor2GDmT25S3fCEuC2/xJW7YDTb5Tct8wsPYjGv7F
TiKpnnZlH9OCIPaNte6v+GjaTzmFnestCie7H7R5mgEKsFhZPi1ZMEa+nkSqBFmI
mwu325dgNk2CB6s2dw6Xzv55QHuo7DCuvBqo0RSkqnZHc3M/TB+TsMQjpMbS1+OW
+2eiCAjt2CCIZj2CcHKK0BH1Ilh0aco1R/TT1SJWVj35zwcEyzG6PbnuVyZ3SVtw
P6VSG04m69+NC4c5N6Iu4pibeTKTfCD5+szWzvk4MtosVmJAc0RzQYKZp5OV5u4N
z3rF18pGlxb/NSGMzBlNxhn8qQuKSK2lD7uon55482mFuF72RfTz5AVHG4SFVRRA
1UgqbCpb7GcSJ0qx0m15AK3PDSIgv4gJ8lza6NnMAfZhBVNjxLwZjPlZ0jGrEfCZ
VG3O3gTWMxJ7EckbW9psRfyUvP24OTyXvElqwk7/PTJMP91UCCk4t5X0FQgFjPsW
QA/7BajDEeglHjdLpqixpAgH4B7/HR9yqXcDEFa9KiQra5No+NJFeDCPOIoL3LFc
4uUgUkWMtbaxbnv2Gd107eVOxzFbjPEfdVxKArxKdX9un7vd9I8606Dj3QnZ8pJX
vkhux4gUOaINHr4cgPu0m3JG5M7meMNyL6d89LuW4susKNU4f73Shuc44QWB4oNq
p44CJLBnQKqdoBhRwkQVWdD9M6iFY3uzjMcccz2E9lGhICyL7qMGnALcjtFcwu1g
oWvCgakdeY17HNTYMXeV0ctSA4dyx+vGMGKzJn9YE/VHy15fCNZbATIheGzyis2t
wMEQna6j+pOmZX3p8HIjb8+EG32VPURd+412dP/lTpQyHZ5mQxT1dPMoSzhuVWy/
0zFKL2XmE9XUDIQyA4b3Pi3E6TMbe0Gld9kBueJRUD6+QptqKXJPb/My3Z6LI3Af
YWpGF2j0z0SLtZjkGLCG+HmloHKuIw/uWXsPcKdTdb9Q4oja901udihiHyUF+iRq
Wg9jCDY1DfYeOOSMLpTLYP/emI1/XwLMjAQ8jPPGsZPkSZojbh5zIholG6QfSpEo
Uz6sxHTd+B2hzS/qFFIZKwdVcovSfRUQ/cQ7nV8q8Y9PYIjnOAmUOlxzGj8m+vNC
HUap8rXJcfeE/8XhtObhOYPqPui+a07P87EX9+AX9Xl9T1pgtqm3ww+QdLKkbCov
etc8Ke/Q0zW8sKZhllUZYEfMJLe6miFTUrIFz+RN77lulrmP/YC+LW9ahAHwTBSx
dU/j59Db3fMINWb0LNP7l6dSmDNUnSbOjpEMtqWNOt1XI8cKu/dWRqRQXe+mCdlj
Ua3kTBp1BlXhNVPeYlC9SYl5nMUJSgSF34QRE6C2MU8mGmn4QOiF8PELgTaYA3ex
VbEtQxVV7Z67iHcZffSR1livEXsIFxDxU8iJrESqxdu/hygNDwWAGaTg1xOdkRrr
BJHWlF1HbJf59GkRHbZcoCk2ja9drxL+tEjqwJ/JhoLVyLMYaGX4RnIssKHVATXM
sGQj8rqPqmjI6P2F7QwVlGiyWh04u0mjJiBSbDSEYRLJlOiFYGhko+zVfu8LJZwV
DUy7/kb83NdMqN0QqsZICMMzbXy0vUcLA4e0UREbDiVE7CrlNedgT5SpM+YqDS6q
BQ73Z8gOtI06tF87qOUkHJGk3Z+2r4eHyNW0zntW087LLgjYVDbie5y8/vd3oRb5
6JLxOYq+yoAYn5ndV3+f3nVNAsM7Tm5d4uNk/k2lfeDRqJm25gnN4FXf4EUh158E
9ihYF3nmJwgDQCJk8lkh9emvpBIZi6OLbG3bDqhm9EcyFv5El/BegAx5Sli15pl9
+rfPypUMk1r1WPZL/Fz5srI0H0LO9kXnpSdkWH+GryhDG+/QeLWT1cj1wDmimRJx
vPUoJi13Vf7S3NLFS9IizoRoeGdfG3iOLCJmLVOitJqxazJGp3SpulczHA4UvdFX
DTpiGa5I9MIBxqx9Iy/o+ufJ6Ksf0BLTJBdDDkhJ8+Vzw4KLAk6Wn1yOtsokq6Ze
Y8Je2d/iDYYfQigTRQ15KNqV523QahJskqP8pgheffUpSllQ1RbXAdHaSlgchVER
netKnMEocwTZ7JKWLOEj/FMJBCNHxiOvPFxqUcKhUp8ekzO4h70bTWjjvD73og+j
WxYWcv49Cg8Vhxlo4PhoH1TOJ0AbnlWzg/WXLMdc1Dn6NNNoNtSrWTUDWfogCGoD
3Vi5F4GLnXmJkPYspCuC+11RdSvEYajfxbNWKuy0vVOww2PZBAMWquYvHlbzac7k
cz2gA4yjS59eU/6eTQisJhw/HaJgKpVrlRKooUqIpA53pr2MhFGYheu3DbXeXEYK
rZti9xhaBu1+x+ZDxp5y+0i4yMa3cbFYM9YN4/KgKnPENJ/5OZHD1/Ps51E45hrX
O8vDPdQljukgfThVVHhJS2NOh3PuQWJj4hprVSHYi6H8gJe023xWXaE758k7Nu/F
+LzWyWnY61LiP7j/rUkdcYGk6fbSr0subKoUXrAKXfWVpZ9a6WIlMVWpieX6P0Rc
mIOmkJEVWVk4AOFDlyfhHX7xzVSryXo6c96DF5Ge6LmDRn9aNpExPs7QPzBES7O2
5SxX10ySgKaL/wE5hDgoe+Ry9+iUS1hmEv+4uuIH6DJ/fEJ+J5M0hopNrrDq1l+a
WBIl1IKvf3A8ZI4F4g/wq4ZeCa1AscEOEyVzUvWAKYbvJDjhSqKXaIVLxSNbKT7n
4+9ces4byLp8IUMo1h0XTezTr1MGiZ91piVuew+s+o6zSat7Xnan82KhDPHNDLV/
d+DJXaqfS0RdMQqliltdpU/GXvMMF28skvx0frYc7tmnMIBUBXTD+SUcHK0pc+cP
wmfzPrtBmz0caSKZmLeO/8uPxAo7WMGcO80VfRh+3f8z4pcmAYHPhlvHczWEMyR8
/nrSjeUXtB1sgSGV5P3ZJcFU5R+SKFFR/jdg2dnulBrY/AvvJTu96vObnudBy40G
i8DDOAiWg7C+o6Hscmn1H7b19bw/kmUyDHYOIkqWJwRf1/kbriyNSnKHHa12IFSW
YJi1KydEdZgfaJzNtA80yHrgfu5LGDmnIgSNbjLTYZp4Ph4UKVZQpotIQ+vPA4MQ
lTJkGIhC8BsRl/5M3T1pYTcvnxx9s7Ehijjlz+WSobKkVQL0KFK5lPmIJgqSYMft
1EmRQd40YT4f/rnIAuXRlaZ9qFmwWbkqbeq5WAXAC5ByNsjszzN8lv5J35QR67w3
ig07/j5ETrv0wEsNrrWjsbz+JfOdI6IxkmFpXeObZ85kU+fv1E7l5U0CBPj7yAji
G5He4LVokO84DFddVu9CDpVD1qCH+X3AFCVazVIXeUWw2ToS6yfxgk5DqeRvpHmD
VnbLG81oblSdpUkfc0ayo/ZO7KtI3DM1SYoHDSwFvwwXz8MxqQMKjLQEzAu8WADB
Jv8N3A4r02FK8Cx9HoEipQsCOsN26nUowmZx0/YxYs+Y5P9PRwZ2giNbZwtFFgMt
s7fUcPI7SthSHzpc1jsEpj2K/RIJZQh3oNFyGrpGAIKdl6xk/2sMDVWexWjjgtZt
depGp5H67ISRR/eiavQzComhI4hg/5pJeqgfcX/X3V5CSoQwq77vAAQJv5KMV32S
4pPUffWbvw5m1w4eEdDVgD5bLnpzg/6d9z/aU+z4i6KiOA+0T1VFQ7Ue5Ljih09A
OmQ0WrgHkQZhXgDRWBv+zi/qoynSiWx+w+eVfzucDvBU0Rk38caCZzHBBs1yg2Je
aqr3HHeOH8fo/6BMuzvMpvu2J65O/R3UN3UhZgqQ8hXrK21AIbRTE/HFpPgx8WIg
rPRC2L7t1HM7grs3hyeCWQKEfZTmhwrC7WNpNh34sibx5UPtsb/09/cCSxSt37xz
ZexVWWkcOGplBMLj50P2BDSMQ62F9Dq3HtGMaOYg0Q/1FsHNpGtWe5UA1uwcscXz
3v0DqyTIb/KFU/yXe4WAI03E5uoBMhQ0YiXGQLs78cBuA2vMjnMze9n5XS88LUhe
mJ30YgbjNBrWEP0+68lBN1xAk9gjFcEIYtmstLT8b858c5z2BlEQyCWIxjkOdAA5
X8Prk1rb/GSKOBztTAkEx7CJw0xNQ3VXE/OuATPtthXI7vCu7tWglxJQl9TskbMb
vwj+CfypBKt5btxCqCbNXUxxA2trK97OxozJP6RckNsWLPs5eWufMSimLbOAv49z
mSqcoP6CpecPDyqdiVTFMkw11Y/AwJCE+q8g+L9IW0NzSnmFfoQsHDjUowATdhRZ
hjaV4eaWkR2jkYB8zm5lmfCyGpG4OJ7M5OUGPi9b5dljIjIwS8Q2q/Rktq84I0Ru
Soaz++ejtEz0vF+87HTaZtun0icFPGOL1EIXSfnqLXOJyNQXgv3LPheIW82PJAzj
AErqX3QVXKwK4FO/jIKc5S2Pn6+Tg2ktSf+aBBwissW0BHtWEMeF9urW0B30wRDz
JmXQCHCoUGCKUwPBzWVNpxPAF+yqFmRqTZ34e4BY7j6o0YtjD9ShJbsf7+IfNPym
jCVHoO/BkuZkc3/2OaYq28ezwiMinFVxz9fVz037eTNTFJ6+UuGl0Za5bB6VrDqa
YTrn7Rele7+K9ZTXTPd608TjBpN658KbbG6rrfrwCHg33eFP7Nc+Aa5pIbMx/B65
jSO1A722jbjaVRxA3VcnmWqy+Nx8NC95/c1nj4FzFM+HvObQA+78UftcDwg/gkRC
/XhJ0/9O4mr4m9VjUx0ZR6TM8I2lbcQcKIKe7spD0Aie8BimorItN3Sp6wTDaiNb
blSTp5I6oYWmNFTTWzmxXBt+T5TmCo49ymNUDq8GsGiRifrtMXGJcGyllkt1YMET
dvIKEfbq9A2ChRh22kMoyGLulxJ8BRMMUjbU+g++iYAaBVDXNHnjudmWYplaZ8uQ
0Mt38RBzr2OZPw7KJmeALRPpf1yT7k9uLdjvySNvz9yFV+ySqKVAwPy4NeVyRxBj
apQSetcsiYEEABBH0GbAQDcNcxTX0hbPo7fFZ9bRRi1gu9oBgyQYLHx6/0UBxSYc
8yZK3ybYDqnsIZlkwqu16nz/Vsjrc2H6bOdpoPXnH1GlRYq/Z3cyjvnSSE6Ks5QY
PRTWfdllW4v7Xo+Hr5oVKIIAZ7MCb8YE50h+eTU5VOi8QYoN3G6oioDbZMLs5IOT
IImLGL6o932/IxpJILKGQiTYNMLs0m6UB6VOGGk1bTNuRk0t6YSZ0nVRYSr1J62U
zC8LCIkr7UkD3atkZbVblV+rflqejgWQM93ozidEdIdTP3u93BYtmBBQmXB9FBZw
NsxEhO/t+/jmVIJWkmQ7OLEgsZ7phj2mOWgQ5WWMrthnzsoRXUsdu97brSUQRG9a
vPYqYopHTNhI/YEJs1XtSZNCjJfcyJ7EQnkINCbAkQPmPViJVsiWLnRZml/xsm/L
zXvAQ1L+FYf11s37anINvdS7cmbDV11Dp4Llkx99kB0HtrrUQGApUWxvK1ycgKXb
pKYh+G5z1I5n/RV4B1KgcVXVOY6khietVuTH1CjhajFAX3EOYu59MzJ9BEj63KRd
lY3T2K9B4uZvG6Co5NKx/lqDymPDPwR2j9VQhurEzm5dP+J7pRCvzI0D1p2WbakD
pjBqv7XBiIkCU3w9hDkle/Yy7aGGvGiNAIm4xHkvyX4IjcTYiBxaTBGiIFHXppdw
MY5LL+3mBMNa7+r48XTvhjrDaThBOjhmPhtOt1rD/Fyz/aXhN2/TUTapmLkw/x0R
8W/QlYnQqYftocRUrgtPG9USR2PFBuCACMYSOp1Pe19viXZJi9HPIKtXxpHecHJV
0HC7YoJ3xXLV8g8QSEyAHxzDX742/jNEmtdYXwegu0hUKo7KSdPjIjKZ6AcuH0jd
gFiyDVkbdAOBu+KDFeVj7hC9mpo8xce0AogNM7dKNZhoMkn4fGXxR2mbkaSJNzMs
Whb/4DXSKJqSoPH4G+0ehTjm3F+aPmKZKxJvytVPkfQ9Aw1xcazpyvF+pgYOWo2X
dRjRo4TFHVPUEZ2GyQHoCtCJx8qg3sGcVundOb/X7SRyDU6JN5j2j9Sb/n+9iLTy
5c3C61cP0X/d9icXL+p7//FTsSsl8CnquWO85dmWVir605b9KD86ESztqjuFSWhX
z4qUiHSKYvTGSy3iPQowQGF7Dy0TuNkKbQEQ+a/8bK1a3GNtk4nYK5etRmxCmLj2
gH/Rmwa/jmEZLeNyjzcT0Wouj+6aYlCSmHz9mror4smu5fN7E0KTWC0kfCwEQOT4
YMHG+Qg/0PjqZx2ROwEKqMmqOPICceFXqDWzCAtgpAXL9czpuuM7laUcnGIOV/79
uvkYu+UXo5OjE7gff93X2iJ8kXtYDm8XEiOE2EBUtosP16cFQNc8KQ448dejRubS
FvttetAFZVHbbCC4ikC4KujTkLJjpxW4z9ky+fO/L5G+tCLyAT6qThc2AFy2UCVK
2FUzTjKnaLSbdkv8w0MS3tQNE4PmlsjrhJcWozlGTqQsCKmkPs1W3HPsq7gcd4mn
i8PtWdMMaMwrjlFz9AmDf/xkRO1VsKKuNHA23+V4xOMapFpi6bH7EznhJxN1esuC
0QRe1VKmGg/LLX3uoUqQsbRkyq93wX2e14RErigaj461l+xcugbhu1gtFTWEDyQv
hQwi/MOL68D16RC86thLQrIMiDrUxXJ1AS+DuVfPub1rdhYRtaiuGo1nXNGEC05u
4Uw8x31JoT09iaIISebkMDHkja4Tv2Pqbe4C5y5XvX4z25E9iEH/EAfuUaOqzIcb
GPPr/vOG07GxRneKGMA5/R/ivrJLSuMI6zFu/E9x1PkUGvAdvjanExBD5Ur9bt8z
/Tcg7E4LDpu7hm/4yDK8Mfd7YI+5+nOKTr5wU4DgAIP8gFaTxPLW0m0UfJwDI7jg
zv++TVn6lkZH5MO9BFL1ivERR92cxq7+xnlJbIIPQM440RmEpu+bhGxb3Flop8KH
FYyuHndSWyXBGVQs5dPoWJmioJb0p/6bBWUqONC7sBCsr9LYhefdwi63uD8JSxId
VfaU23HqV+hMDBaeWJC3EBijW+/TqIVmS8FpuvM8vzTqDitGH14pGVs2Fr4KjEVK
mcL5NjKuOLskk5tTga4cyl+B+w97auep027YDLaCAyzqsP2igKGiL9dUlswviS9O
6ya2nN68kJelMfJrqY+4UXB288FJNNE9/mrm/g6yjO3OSQnKbKDE19sRrodDOcvG
y99cwgXMR8lpud72To6Tvjx1pehkHASCrs32A07V62m7+3me9nT2BPCI9He0suVv
FeP08x14XBXXtlOVaRrw4wvZX8F6shhAQDIQpcvG/a7HMuqFSpLnpFvQuBZwaw92
ys0Jd+K6qPSeEflBNDD3UR3OKunX00F+jsfdE6QQaFT3gj+Tm1k1r1n4pouuQm97
QLiCbBefvWGESi1iR/pVbOXxoEleBm0k4KAeIocSw/zeqieDFnVpFdSaeZzjewew
b64TxS2gdWGbssFDQf2VhobsKWUYsFRq49+ZgcNdiD8+6NMJh/5eJ3lXV8sPjhXp
7u3s7umvMjGo7FNpITLlyFL/HUDr9fDVg9Hgm0aMBuJgVpr+rOIG5QRAGsLelD88
U+dplbfb8FrI1x9AigO0UlCc+CYPCB3pJNYvrytVKvqB9bHYt851yC94cavSnrOG
X7scruge8T/dV8UtlO/7wuX2RyyNgNhkz3T1vBHV8rKaCGEcxxTwXVXxZz4SDp/S
AfS3YpMmkjTlgOM+PTtAFE+E8HnX/Q0CC12igpuUyjrEJh24nZxGMoLtjo/p0GLs
TvGQGL+4Orgj/Yk7X6oZHBiNnWiZAzQdrRk20iKincjBL9D8Q2LE/r+mxhJxkoK+
4g+Hou8euAMYJREVWmd/JBosLsrtB2t57GLUaQSdm5JqMbcKZGhN8+JokQWfeepC
iaIwrh4QRrkjVLsIGdp5uG77sEnkQ2VQ87A8ZPN98/x+KH5SCtiRZCWZ7RhZbWYf
fnGDBN0+pHQY55ZwqhPAI8qYNc0dYoeyGvqeZaeZ/zmhgdTDnshTEF98jCskGtsa
iCydvRGsNKtRHbIWAfM0pL5djW/g/Kot7eY0vjFPnhxwnUENBGwL2q+m01ianuP6
vFdDuxti14Hq9HoWGLHvO8N6qTqiCAio2EzGXw1N12FLVadwdnsXbT4dhydCuv9h
ojhpaga508DbzXhgqIyPC4Ye5FxgdHHo9Z0gJG/6+jnDld4lqWHk6JysIu03C8el
pNqKvK5qQAmx+xb9IGeigrEyOZjPqJpQMw+hsVtlPGacTqLMsxDABuBdE9MetlH3
zWGlVTutS59PX2X+UeE4HjXBfWuQyFkdS49V582PNsk1G72JsE+I89pa8g9//dlf
mr7r+5mcSNkow64FQDV+BGGbt5NkobqjXNmBm6J0wcxcLZmGEOGkJDJftr5KZNFF
7h0jI6PL/bKrkIxDrHcatVQK5phGXNgqJpeDfdq81P/0hfgd3fFxT2dhgiyjZz7x
sE+ag11q2LtrUQMbVdFvo//ZuOgcDY0sELaga2m0322uxjP6TeABxmboSSgx2NLE
mwuXVZekFubQawndI52EFzpajDCBpv1efDtmerzEcEt+DXRKB+DPuriog4XFcys8
8raMga1DvCE9hmRF9u+hbZcWazj8TF9JxnAKRg50m58RnY+MjU4R8gMX1IW0hKCR
5g43CtiZDovMMFs/TdRbHN3DNmpYBf+S8Btt8P4crEHhIx0/zDvS1IYccAVdnqhC
3TN+AifQw0Y8aBcMWyZW0ccGmnf3godOm4RNiPpVZ9rKRdVhihUXveWhuuOb5ywV
ySEgmUDqTwQg+TskETZW48YN7TByUxBoPCSgn78haginM2PTQioHK9UJ4hZIO294
W8OICeQepd2yATT2Ca0dhlEkIS/xkWl+JIc0wbMORo+0lC04NYPKkG8XFmk/Ie7Z
cwc2I6aZp7//66ZMvZyXbMeeAkzhcLqItJmyYk3k4bqZp709De55xzIPwigtAqkQ
9gkjoUIgtH5I2Whz4eeSGmoUBir/HGZzT/GwEY0RC8bhEvXQ6nXZWbVDAZSijDb9
m7v6pTb0USXS22kc+CkXkYeoYsKiIHtZfVQnX8o3kc+wSfMjdYVhn21j9A3ykPkx
l7njkcWTSGsPZM/MFqq4pxIl9nju9cOk1h3lw0QGBtjCMxgx7A3/1udKTxHOx5cH
KPbQctWVJCl2zWem1S4nl5azf9JeYPNU+KLvlU9vBRUOKcaw3aX/eu7zdceehSkY
3BdlhTxjbEFn4zj/Tvuii4HxXHYQogSS3wBdJi0e7CjFvcism9Pp0G5TFuyV6UoW
1QcnD45BC5KrKxFQdy3trYPh3Y0wNvJlpk/HqoF2bjqI2pyoOIYiws0tRs+5dNby
MbldTt9r+n1bd/RnBl6aS5OhStmtnhGIUMv/XeRRnRK0c8S4DYCaWh2A6CpFuvC9
ebCM7Vb3sHzsQ33EQS5A5PX1Vk6z56Bv9VVzJ/nskwaMg9hWBElRdOYQHhkhdAWB
HbDb3LXCDcAgNTyzKrU97qzTMdzfXNnh34oc+QN2hjbefWOHsfnf5Vs0xlJDXxab
ebUKS5sSisbHfh8P+aihm3RZpw5JuYB9QrLVXJA5QazMTEMSBwdDSA906jzJDadg
W2mEt1HYGwP0wi2uxzJxTimR5tphULL8sIitXNyplSLd6XQrXVwlLguwLuDrTOK9
j9w7Qci2njOhiys3iZqCEnVwOaK0KPndUrgNmYwz+ViA8UnE8qz7G49vdVFa4uSk
EctvHoBlIaKPSigeNqazzXkxEnF1lQZUcRs/CpnXsj7+2QJvuUF9CAl8nxnVIGxI
vqjxJQi4tP3y5NpRhg9qMitgjP0xHAEbMnUWB2+7GrVYw4/4Wgy5Kkp2C4ZbyYOS
QOWV7uq5EF7fqs205rO/WTQ7HJpARNBVWuX1/7ZWV4XnfS/EAfVeqW/mSdDkd9e7
82yqEcCEWDn5Dmynz9lYUD57m5n3xbD0M/9o9vrBu9wLED9rnWYejVTehP+M2Y9H
3ZO42mWIk04ka8AVYXboEDDZS36IGl12iZqidqqEuuD5Ggicfv4o+lAsAgMjMJQt
BHFIpHdmS/RZ46qKzbjIT/Wm7v51OvHsXHNstRPABJ3HHOFu57DJr3Vm+33SnrE3
3GQ5TB+5Ic1IhCJaiKFOMU7vfVMgneTTTSN47v6e+QzjAF9TZwvlD26Sf/64gxdi
OuXvcZIhfN6ad+fwPcCCztyJdoKpDZRq+9++PN5nWs9T2XtXzcWdj7bpnprj9OqJ
u/I51BeIsMmbRTwJPSS67WemQhimWUF85OPK9I1R1PXMz795/NeSgb3bCkthJbQc
LK5rCakVWulBd7iSzAoViwxZDlgd+CvrYqiPOgn2t+AmYVv9uDpRc6w4mIbmwkff
GbR9fpRQayfL5XrtCTMe26ZIPAopuXUOLDyS+D90qCARqQqyklTh/JNs/F9v1/lS
bCd7+DlPgqKniItz5LoLU7qTp65MvNnTVVDtZTpU8763FPv9vF5VdCNIhKECEIij
9CfGvJDTqc2ayiwvaIb50y/oSEOYdZhGbdgGq6gPRku2lbHRuEKb4cqukIH+5dYq
CRVGoJC27zr1juFp3GYyHaCsSCd2xH7FeYaYIO6DXEqdiOFlI9kMr8TDJCQg/4zO
2M3C24RdGfn3eO0d3bQmeeWYBoT8f/YEDAg/qIOTRTe+c6u7kAaHs3QyhurjpQDS
YHvwVwtT69UAovjS5xVmzMkw9ZsXKbJtCDf2ECxruro9IihhTkX33TPYEX64BQQU
vBQ/qtZzL2+1LM/8kCMcB09Ab2tGqqf44p6bM4zwMakY4ZXUy/HwkQcFwAd2eIYH
guPKlpHs8hWXjpa9UKotgYXUfDsXRgQW8jNqFIaD84rQxtWPL96FVbjr2T+8oZOU
+lyFRY9HDdfEjAE9jOXcq2JrL5dRclIyTa9qXoTZjT7wh6Py4ITWJMGC2bzAXCg1
Je7fDBVBKmDHcAbhsfCNrCpAliKhIBMF1/KIoe2hrcDLWlRwqYvRYfRwGBk+k1CF
kM0PC8ycT6sUEyh2ErfvuhYObVwNJrINYKmKwMFNPW86ZBViM/F0kx1NfLWVte27
ZzfLQs71n4tkPCVvNz/EwQO2ivWZGMqZHT8qSlEMJjuWVVzV9y1TyZH+JmMyQQY+
CGAWuviOjXXpZFcZsu8vQqZ/WhWQLe1b6fNKdS2yEYiDpu0nvDTN8M+W/ZId6BMb
ct6/ikr94OVz6QmaexBkEB6dWSjVxFXi+Pd/LBwrxpL1Jfrb1Uvj47+12XTI+AYX
YLkpr970CRhIZGVYAnrRbKQwjY04rq9LhW+pC4zIBQoGvtlc8kDdZJ4so9jZVW5p
edxvoQ3dXtwRBsgPrq3ygOkyritlP5z/Sc84KDsi0v/OmYV0z52Neo2PRY9ygNyp
schdM58l/QX9n5zpcXbQ+kknJqIH5GA9t+XxHOZ5UJZVssiJnbyfomTtvGQ+tsTE
QfDHuROcjy82G1B8vQBOC0v3phTHzKPl4OYugwNpP+uS2HvobaWmAGm+iQquMtyq
NQU5NNegFNn00TDnei4c65yZTGJzHLeU8ErT3uiYXa0YAmGT2C2DsC6IKRWihCqg
IV9ViAPG5cNqeNXHbkMxKsl5HRegikEEgMJ3Ay4OP9mq6RsiaSKOW9QtqKtUMLsu
wJNxAiOTkGjGaniRLNFJn+72emDI4H+SSRMAfEtNnjpUd/ShflAcJau62lUq9m0E
zXPP89njYntTKyAUwkvv8pt2MQfHn872w4bipRO8RBCK3wZx9RQ0+tUdHLN/S7k+
Ca8wAoe8ek7+uRgBjbS+GDWpjen5vrmYYYWKQvJaQlEjods32I78BoHlyRUfWqCt
70hMn/PvW+IDi+swedtDHVV9P3xbz0AarS24MLp2owasyLcCuhQvYsGr/tDvG1pM
fmIGp1/e8HWAQqVjj7cKTixZGYenvMGWil9s9m5JJmc25/pbs+bEvkrhP73e8iV5
Yahp1PVrLjhsLimlfiOtIDxGqVTnLnJaxgir5lUre4zQCGSYAjqW2SAYR/ht00SI
xPrBqdVZ57BIjHaeC+SwBbsxWNavX19w8M/laBfPEjWB16XOr+zMJ/HPwVpXCUo2
yOzivfrF//1eOZ4SCNWqRMHzmaKCStMJCAsFKA5dcAP1awg7jFRLtJw7Ge35FlB9
tzoFoWyvXJxxK/J3lz34UnezZxEJn0dTRpzJKStKJgi0S4MV0CMqpFVmYiBdTbbO
F9jr0cXbosMPLCw3B0Wdl0dQjaBYvBOsep2Va1rto0Pqa23QJBSM6ea1i1rcluE4
zVMMuMoDS1fY4Nx5qyWebtuo704N8bIBw0Nj+WcGiYWdu0R7YTwnM2OaH0RYpZ1e
klg+crpNquPEo0L7VRahE3yQtui0Cp45RSM9J1kzVzxp3FACBfN7PZHw/C5/YCr7
Y8daLfwaWqAByxmPLr7fiX/HKVgmj3ytWnNRNguOZgi6NrBHP9J3tfOW8q5PcFu5
r6w6EbrB7KFTEl4wqffcAavO+j1lLxA63oIrr+PFZN55v/Q79Iri5EORjmDgvNln
0Fx7aaHofk0bq3Z7iIxAALgNrYY7/WeSpTvfam3kBexn59Vw0UpUIQs8PdX/fobw
15UEeuIzOwL45ZYDGupoKE5iAxNQnCd1sD/qfl1Cral93IvvfsREvsST19BhP3hq
PMzw+H78wyLxCEHQeZOzSWrnJ7tlgtmKtlLhTJ+zOCMMdAlMCKR62I5F/hje04Ec
CoR+0hNSAFLQ2gIFbexpvWnGg1zCgJwNigMaWq3UFQZ4ZHM09uD+rCU93ePHqa7a
Ke37riWTq3sC9kqAfwkafYLCAEqCqnYW8INtrBwWI2dvPojZTbmAcD6HjhHUwR7R
G8Zawb8FNqaC2geY3/5v4Onml9XdLF9usKhb7iJW3craJMNECaLfCDRu8/YrDLIj
hZA32vxuzDksUhIdI8QlYfWidbDtdROyMBRDRVn2YYfUneewYul+LijQoSf/KgSh
ns8m0Gl9NGKtTAYTNf6PgBs5N9g+qzhhXf+ismLNc06mHOdnzDnbaIqwlHVrSDLt
1aukYTvflhioyL9Z78dOXNvSOc8zEhJzfHjPiO7SPCswJzRTUQeAUn7jRyWxNogT
rbgYF589dP8HYVvJs/bSdpnI1iedAzBbQq3qZiTootqIPTwFm8f5dWVPXzbJ/WJW
Ur7by95tKo04WACe+U9maMhec3S6CJGD7b+S9RwnR0to5R+pIP+RIXgPFwTa6XKV
VQwCtJ5gq3BBOds0IC1qovksKaXzQkQYrW6GyKITbhHXVz21bQtl/O1B1HQyYz/D
OhgGB7yfzxqQkE1fxTGEu/N7M77MCSx1vxzEdWCHB5NCI69RqAEoCjFfu5SI3xyB
gOmS3AeU4bruz7vgNgsk0UxZ84UOSq9W5CuQZauz6+IxT+caIQaCzw0YovCFdb2m
QU0VPSqlF8yq2jKPojf96U6wBmm+wEiZHmeIBqO+LfGYfYF9EDgnOvGCE9TJkkFY
vZlFGzC2D8hFKDCIjuLj06BeFZM3y4TrFU4zPLdem6eD+iQxgtYR6g63/DDA7/6R
pIa4SCZDYFx27k3xDBJ4/d759jXtG7C/UwhUKXJqWsjzGzHpLuVPZ6oiwbMbAY5T
g18A1+Eq4Wd19mXklZzmJjVi3Jb52o5AeFHC1Z/QweDxI0am5hVDfRJc1rR66R/J
knKreaZw4Cp+UzANExE0Rd/XWDtGICzmOPKOQ7Vvz+g6xP/NQjcK3ywbJ4n9IAV8
3bMmtCryr5KxUiAg5Dh2KwU2BIrXAuk6o654NcZCPkYldWqr7x7UPG2se4+OIxy0
/zOfuG+2k+ckVc62/nwwpEi1N2x2eUnSAXYVIG7fq1GTRHVWfhK0KYxQCSzs+8Mr
1giVP3RwLiuF7CVO6zhz2zMf3Ks9QssIt/QjalRsjXcfeNRbrzaw7NUIu/KbuTNC
2yNlD/6o8atCLicVKlGZGkTzHa9M3ta2yC5459pur7OSr0QWbQNdNl8aUt0z3In3
69jVOr7N7yq1gZg2Dpu/YkG1TZ745ypaosBle3AMFVDY4moiaUSAq+7KaAPfP1AY
Dx/Jxe0ovW5EVziLN3p3b+i2Q9I3vYHnNwF2xFb+SkZMW/c8TZ6yj32piqqu92nu
BW59b9sUgwyRaihA2UBkxnLoLigzyYjxZQXQCmMURcY41LR0UEGTwmcB7oRh6JUP
mZEclolbHMse0Hf9ZcPIHlibaVUqpA9xhg6zG1QXjUYEqnBEbF10e5YiiuTgZTgI
vX/JAmlMiY5T0V/P9Ymw6o51y4gfSRIRUwWUyQ+CdUISYIhl81ktq3fwlt7VUFuS
x8YRiFZtQ1hs9exePAphjR4VpeTos1Ng4Nl6tj51rJ0kJavdYsSpJe5Wy1Djx3XX
OC6iTHamzsTqx4hNQ0fR7daqOBMfYvHjwPI2g7JdQa8j5WAPrpt8iolYD21NBNL0
lK8dhn1cgvja1Xr2szuDgXo+Edlun2R27k1dpmuwC8JX6a2ati5JBp4Epec7BF6G
M6KTRGU7UnfUjNF4w9wUxRPBVX2HTACrzPwgJNOp9PMtihL4f5xU3/CzZD+lThAW
0tw1c0s0mouFGWw/gnCGgUL4mCO9gbQ9eJojk4PaiyIEHVTDolyEIx8gBrhO7j6+
ASFBwlZJcNrgIVR5zMwmJ4MH70W46q87yZ+r56xjuaZKZmuhIXgIoAvI2quFiLiS
x4nICYqHSBhYKRe88brXh6y64S+1eW985sW24uAj2NfjKJGKAs0SYj6Zhp6RMLbQ
kIakzRD+t5g9u99jiwIOPczuwe3CkP51Q1ySXUDkOsN6o7q6qcx+VFrwE38HZLi0
EC4AogkqyEttEQADlh+W9NmRGr7MBnnfMRQPMe7jOdPp+9pak9qopzud0JTTcvYM
KuOWgPhbWztnDe7NoQrrA2bGXWK8Nt6xhYkg94aXnTUClG/ez3X3UIVWfo23TRYx
GZNMp5ggeh3c33JdIIhQMN83YkQE0HEn7jLcJf5Eu714HW4uYxa7mUS+NixQ6qZL
NFABiT4y1MSWjTUMAZY9iQyYtt/f02p3oEFQPP0uLLFbSvGOXMOLXAHFtSZX900Q
h+2ffqgv1SOelmPsolMaYdmQbbVwrLXY23CECSxKJl3ZtTMzVYsDvqq9/bahooUj
R+tjjxi+IZUfDVsxRmZLK6Jx91e109gJhUFH4oI1bFNFXzu85Wb1FnPgIzKq9H38
sQNW+BHUcZca99Zgxsy7cKTcnyAXPBZGYGmWws5OdYqh8SrFfnmWEZmkbDf9yx7K
tF1q/4hcxnTasK1JOzCuYzrfYfy8sBZ0aMOufSOhAv6I4+h/3NgTCKepSUVbO2Uo
DOGPXa9R5roQU0SB/kPhb1BPjvxdPbufB6EZggc3q+zooTt2saxhFZ4CHeQLeKMD
gVnIsqlH+a5pgzK9M821kQcaSu2GrPcuE3whR4G+DH1yPv0Uaem0kMMlOcdhEZAr
zUI86y8ocdPE0xY4FYMEDOjB2tv7NlTRGTVVkH5vaXWD8tPp2s3NVw3WRISyL4N2
jZx0+m2At+frpWkFuLJp64zCx7YcpWCsed5GewwsiKHqk8JbB+rsIMctc28lywlK
19eSYTMi/KaMVnh9vBNsyCNfvbke0ViyErTIyehDUxIrzj7uqDc9oK8Wl3INtyWM
9gckAff0EuBxvYV8QnSHL+eFB0HtCgTGJjPTZOIQgYMvs/7TUTEOdgKsnvi5weLv
oM6neNwv0rjQ2q9xmqr6cG9zDMHYunQeP7YpDuS+WZHdWoC3taanXfbFy7t4WOoY
AQATr+IQLpNR8OMZvldBkJv6L7Opz9pPTu9RW7kCc6gPzZzUmxRwNYtqMD+Cq6qZ
OHms76cAHHnwqjOPDkWRrZSpNHENAFWxcVztnuOtw1giEV++A+aep2oRuEjjTt/G
z+ICtltgACmiMZ3TOiMijtqABhXoHiNM5lUpe9BD4/9SPRWcX0/mQ93eXNlHeB8x
3NatazqaY/pv9G/7vNKEHyn1jg0Lst8r58K+rkW7Tl5L7NLbrlPc7x62QaE2G7db
OpiZ2DG7OfvKKf4gZUxyKdnUhMz8e7YYysoREVPMD+2C3tBcnnfMYZNmOR3c5OSG
MRiAy/sh973gxgO97dxYR44p75qvK3c/rgGnx33Zvmpq4X0YsmHV10Du9SxkG58s
5FBzOaasqtCv4Fm1RAExO4MLf8Zr+8L6NsM8GvIrrQcqMRKrgnQ97chpG+r2j7tr
AMG7IHhzcF+CtYX4U/cmHOy5TCofEttLjJ+En7BC80dnu00gvVBP4P2W4h4nDJ74
hywqioBwJTesXfdC1vHv8pj2a5vnMvBz3gHw0FNLgZQ7LK/56k1hgzsu4lsjkFOR
Mfms8imrUL4hIjJM15tMv+hbShAoilDd6cnDC3hcEZxh06mujaj9jBso7myBLfu4
1amKRjO46L1zn78bF6vw6vWxzMUZX87QA9RN1TeGJSxMHI0fETS0dxG0qCx4jaZX
nyvfvQjR60QVan8nClPmktdu7t5vu4CubvyVucr+jmBXBlbTXyAe/WQVInIvRlFi
DM3+IH6EVrQmkbaPF0bhCz0MfNZPb0W15hHOIiBLZVxh4LJ/eTtvM5ugvd9qnfKr
LXT+p6nqhnMg/wjzCcifHLgS5AHxfgXGudThqFv2Dup7EZ5X9O0qjNvC82EaEav/
eNJEJh6cNUOBpOLSBSfXSUi8rs1sDg5l+OnIl1vOe8k36BXba3QjOUClxb+viMSS
0u4oWWbHxG6FWW0Ydt/hbQFa4+i2On4pcVmGPhTAjHaQ/1v+CyEqz5+04Rd3yqkj
4QK24Sb4ma7VJXGLLHd3nxPlnHxPkeu3WROM4A7+OSTdtCpYEoHaduq7iu+RsCE/
gERP0KooctGtTlYP78ZAWt5i8411UwjohS9NT8z5D1T7ekGkWCuTlRkC27sBmmXO
NTUH3adE1fd3+EX2vge6+x9GJ/OK7lKAkztorUhS34D26tEBBYzPvLi7IN2MlMXL
Er3in+ev2nzV4FNsi2mP0YoGw9KImF1/jw7drll1BAYtcrLvKSO5oHgRc5Ns2FCM
AsIajuRBvIgiZ3dZkdGJbph9lkataMexHbmZHEJzpxrD/WWx6ygCxBFnlqSlSCYm
wBZdCgzVkjNd7SGIXKQEwef8QoVmeOJxLrcBdwDX2/hbipa2+6gYJh4T0UEUI/80
qneQKGvLDuaH3koPXpwGA9epOcb7e5OQ3m1F42AJsyeZ8zgaji2S8Zz0BzxG2OMr
WTaGt6Of2nubrtB2qpNOq1/05TKbHF/Vkeg9gFn2ex6L9WLxtRQKjK0GnZjU3L2V
dolmypk4Tu7KDclv1EVkpGa1YMY8XaxD0faVqA0I8LEpTYX68Sz46tk24WZDYVQN
Hn++9jXdlPkMz+aVDySQhDpvu1+4nYnbELcQd9oqLIZDKo8N29HkmvYZdIL2xETN
mKzSn/u3jWKrf4WhRUuFbhyemjmJr382lzgoR7pul7tlD2TSpstYCIBousdt6bOL
T+okieG2r2BtD8AotMFsGl4oGHqjyEIJgU+yGjNWCskuCQG0vTWFpx7AQqVXQscg
vxBuxZJX6n/Z4yI+67hB15AD0br6J5uxzIE3AJI/1o3QVgQVjbO5TDi6hNmxEhAo
3XewKG40hY28P9G8COrMJzFMiPeQdH4Cqq/E5BI/VGeqX5jcX0DKu73j34qJyRbj
dLCq9u5Peux1ZPCPvyVVLhl7kWoQ7K+f4A8WidZS0CvgzKgdvWyw2b0XeDEmwEiD
CcFrgguMHr4bZRMFWtwQd8xt/EIhjTPMLUPLDsgESy412P0khR13VwJGldDDHUtk
YCjAWkRpP3/TA1MbXWKjEtERbK3NU0qDJxBcC7UmhEWcwBA1CKhYQ/RSwseCkxrs
o9vguGEznQTVAHpiVyEr8E9WG4AtBxHra/NC15QTL0gPBpzcUnJl2zzc015ONq61
KbUto3UStivIzJPk4K/JEIJEFiQkeLE7XxyiuXiNluOU0DfbDZ7CBCPIpd3ijxAb
+Mqjyif0I6mEPlT5Fs3OeQFXRp28Nj+9a6mycxdVIoWIVhPZ6rW9bK+e+5f8HqAv
7CRhmrin+WKiIflyt8cZy9WvQ7EBYc+kh2FwRuTZ8vaQomt25QLgbaoD18u/lmhq
MTOarP0TtHre5Gna/Sf29APmMvdn7g/lTznB5B/GUbUlmTqEya24q9ChLXL+rbEW
gukwF3YXsFbtyJkQOku7iaDB5xrF+tIM8nDcxLPDhCln4Q5dcuHdlLLRHYs2L7cA
SDdZMO++HJDKtoFqkamYDUuG6WVoE8ZeqL+s5PF7IysYO2g++rJZcbBbWTOLlYB1
gheBntzGOK/t7t4M4Is6Z4n9rDkVCCwnEyG9M5v+4t5YfVSx1nU2OjNxHutGSD52
nqlAS4fu+cM9acwK6QmYOrHZLnW46g95mG4qNwEAYY/urnTrTagMy1WE/3cZIM5D
XX8dvLM/eD038AbM+l9AIL1dfObnTjClUvQCY954rrBA1eNPYStYtwWdE30xCcpe
njqNLlX5xI4Mqy/nfMs1XCwSRdx4rGZON5oTzJVr6l2vXE9XcR0nGGmNrrJ/NgTT
2NykwwO8wJaQb4zcwHNju8+djNy2/VGr4AZg8EVFxW9FAS/aYtySE2c1wxTSNMvg
yL7rG4U/9ekiRGF1kxHYFmxmTVM7p6e1Z4QokfiJe58WqmT6tfH2Xl7McDXn/55N
Fq5eC4q1WlHqTeyl2/oI93iIh6avMCGdhSHuIhq85e6i2yNh1fSTzGP3imksUA1e
0fGZ+36xPBzUzZhxIvSnlZC4opSCVJtBb9YDRuso8Wxt1DbuJs5yhuKPJCG0fIJN
1mVZx4e4uiN5qhI9LSVbM1nR4P+7sE8Vpc7AyGgNqMXVT+fRRoIth+Gphqa5MXsF
778TtuQXM2GoqJa5lM/q5JHzeXIdxV679Q5NgxbbGPQbF610qwerMz9XTJfYWoy/
O8OFqD3tipdhCL1OqpqXz5cbCyHK8oWCQoSJkEj1eJ4VZloYJFAl1LVrDoqdpSUD
tIjnrzV2fnuKjfzNXkHg/J13M91XSq7qBWAEK++zNuhdzYnvS/g7sHHv8xDt8zY6
9BDpfr0NniQPlDPac1/eBxqJkDF3Czd6BY4RlBhA3xN3EB6wHozdVoxJE+/GXNQV
IzyPErCInDY/6u6jZpRxJ7TncifOF3yZ6fnJ4kMx/YLha4k2ALkPNw6GsQna9xAw
yic51XBeoMiHycciezCtWbUSBvYvMduQMclDhUv3iltwWIP6WVrhbItC2wbLFbwU
huG8yDV1P8BayEzaPORztWn85i29x2dUIUKiIL19yVyawYGkBn0yBWoVI4IA1p1b
ASHosQDJthfOxC1SB3HfWIoJQjEMn36fR2/GyrTo8D1n9v2OD9uIdVfJkKOkQhfc
Z3oTJGXWRhZvxCoKOzk2+w4zofE3D5e3fpAS/ahwEK2saWzlUniKg54Y8Jlr3osp
XcHR4S2P7PHE18SVtiLUUb0R6PeeVb+sPu06RNO9T40qcDvOPF5bq2RwJt8ivXQB
RSBlG9N3n+vktu2YKnBrGUFDSj+SPvWdSk01hRMDcQ2QCSJ7B622q1F51XBsHLku
hWBmA0AFfYl7jrs1HNzyux8T1IZnD6XqEw++FBc+uYy8Xoi5zz25r6qed2fwjx9f
PynyUf9MnjoZabcsCsUFU7sg8b4G7KtyzGyQhN3UPlbIKn3R0ZjrcUQ7c9df5RaJ
o1q5rvOLy1Ifi3rwC4XT/VRRiBOJy87UT0GrHzRBCxZPpeorGKBE5FjMwEYHNAnw
HUtkVgkZGnlh1gS+D4QV8bx23gJAoeaz99LPY3ccVo9skiWXbnFSHk9xnzVVDnmx
9eM1ZaCZG+1b9UijO7kUO3TN6cK+fRs3TMLiP9t9YATFFyCgGZlf+oU0CXOD1/Ll
Ow2CdG4ANTyH99wVxTOaR7qRsLDs9VYPcDcy33gTR6AFkM2ZNht+HVcDYcycz/kB
4ApiM5Y+TBOdANOnGRrmUFbaaC0S9TFoLY/roiC/XcSSX+KfstVWEUTE+JdVieUh
PY1K7scXoPNKSUo5OCX+ei2dITTCoYv78BZoYOnV8VDxVfwh0XiF2L/zG/G3GGCO
eNoJFO7zpjRDx61j5Ohq/0XNXB4oP+4VOCZmAqoQBhH0ADUYH0QK/jQdgMtQv3SQ
mLcgUv6r0Ted2/hVHswZs/EhYkOr2o9V9nSKHbWRgnBbkU5lItPOsH6Z3YvwYazx
+meJZ+GMMFHHeRdX2nbuuR4KA+GoxV4KaDTjLwQLhXjnXu19Pkmcitk3XYWTtk3c
/lcW2MuPe5x9vi4wsdROJrHbJprEMZJi+TKBk6CL0mCE79HjhysMkP/jzZ7IUmoW
dz6rAVrv9DUECZcHkQN59WmSCgmrwpvl+m+deFKUZCps1xQZgSgR56Ai7aTt95g6
1nMCv/2J0IsUVmlO7ybk7yKQ/SAdYdsuqKWdEct2h9ZU+MT/6bN1uCjT7lZf9kP8
E5bG7tqtA8DMcIX7CbaKaZBoDD7DPo0Rool1moM5QZgAC4PGkvz6AwgNcPA/Vq8b
1lg28B2DW8iyZDIqiYvQkTdQ7pmGSQ+Q08dFzxm0sQkyYkGcVXX82bg+NW/2a+F3
n9+TmTeKDDICYGrrAjXaqFAxk5BOXcnWfGOHqs2cxpHN1Ws1a6unrsajhjVRQCyd
tjjM9Z81KB7VFXXoQXkUZuXU9aHUAwbVl/ZSpX9xxSQkm1YT7hHTj+6TmbMw5hHb
H4GhXXzWUHGUmf1fOasb82uRuTjKPlnvQFG6lKS6gVQIAXgOUrmcdPysvF2GhMI6
8E8Pm3bey2NuoFfLvNyMOaTvlwjc99Xq4o/rOsfh5Ltp32lty3HyN1Cfih5PHRGn
yQ1zWrGjDsIIuTiNiEJC0bo2hBXWYGswGfKPoi/FbhW0R28QjfUVo0czPVWyThoF
HDNPt7TV4C921hcy7usb0R9+/rcuC2dPjqzKoodZq1fzqQ8eatRH3FBlvq1/pzdk
WthUmOS/lb+y7OZiA622LZC4pGF/CNXO1Mb65GbPY33LHsGX824tnYYrKrRLnlsD
KAmE4HhrgO3XR0/cFydbFp8NHr4f+HWwXUGlY2Jmp7IvjvJi/4fdyqADqkAta2GS
zbY34ZBZ4iXmQtbXfwIsOIA3Q7q2U8J2QSCFbQkd/O07W45mRxjX8W6cwTu2+oVO
+Iki8YyiZM4AYkdmamScHVgFRhv4S3Nc/VZ3BXSubXLYoNrCPbKscn3Yxndnlw6s
9ekDqfH1+ntV5ZqqLFhAaNAMfgJ0q9H+O1H0SK1YkqFOtigqicaSIFyKax8adyxg
SpBLmAzpKrWi67vuohUJ67evepLSGtpqpsT7EshXq2yf2joz+mi0TYtPWdt54rEB
x2Nv4A9PYYEJ+Cs+/PiCxaYpLutc90m2U/sRY3/0ZehffautvXm8E8s5hFTzYSx+
gGe4La5R9PEWprXlp8JdDem+eJdoxxoALMx9W42bk6LpYMkVcCT5aHBjnyJ1+0Wr
VjLIZjEEQ45EX2xTKYnCc2f3NPV3wnZUydqgw/81P1fGITSemgr60tVhIPx6lkOL
L0TNa9IrP/po4zstGypzNBfpgkByiTeIRUxSNJUAzw9dur1TLW9qfqrFSCQfwO/x
s1MMaJvAWK5openhMZLlgNrp/0n3y3cMohwesXkm5J6k+M/TWsEEZ5r17xZSOCr7
G+//GB4smuUWenGpARI7gKnWFR4r6wXEn1TdEre5rnACPa4eUTMYXQ4B385RueWS
FiOn3S4rL0qGznWllEsdjpS0hja8aLRLY4XABGQTM1QTfYMma4AgOf9aaFmD/IY1
C4y6X6ZG6fS3ge8xo+TryqK97eA8QUfehdSYSOM+bS03mL7kxJXUAxgC35QX0M26
f6eCfeKTheJUVnT+l3eRbDgL+mVZqRE4vaC8W6UiH3n68RWglVerxBc5yX6LYtwn
x8WgRS/eF3LNQvXNPOaRj4xrB09n6TgOA7a5EDtRXgzu++H8h4tGjCGeuQT74kPA
+Md9Yg7lxVQWP3b1ZI6oa2bjQhGVOUQB7iJ+7DJE66s95nzQdxvJTxKqDsinc5Vt
NjH4tD0MIKHO7D0ysN1318sF9PegLZmnGBRDm3NbVyEpY1ecapYQ+qPy3FGtpIPM
Z34wyHGrLVnbN/5UzzL1MEdeTuk5p/G+aHZF69XN8vpClNv3NECZaZexsyeLkWDz
f1RdHNX1OCHYbnqdBK0dbbgl0LIdyMyJWPIZ49GWQaUoa03CGgqqaE6VB39l5enz
5RkCtCzMdFdhyvvYLraT/rFQgbA6X4qvvi3llPAnHk9drgrzHoNm17tJF3yML6Uf
GsxUO0AQMnBZF8BtN5KQX9/ZqdoPs6dQsYeA89IUC8C3zRGK+pMkaNCvIckL5gCJ
yUKRXAOzIZr6sFuaGTGa98q4T0gkCnC3wBmpJUPhAxvNr6aOH4DoK4A3w+SToXGa
ilVCJ60W15WVydFz63btCdJGJ6T3bJbn1J1+tn9FMTPabTlkO+cpSv+F+f2TxMxB
MNhHwLs6eOYFLq9CQMTpSThJQ1benYupzHsd/bW03+9wk8LLeoPYOnwgepIgoBYz
eAvkjARJwsZIkcO/j964246rcnSWnHe3rOhX03f7FuFEY0G29+6VQob8snbV7keS
S5Rdy1uj4/ijibgFnQ236ycRRjx/cTEpLrLbFsiescuKhUwkepUIWhoshdnw1Q0R
XsQ3LwO6Enoj6xoTjEBvP7viNLByXc7udBdn1MCXbsJX3PnZZmwvgjJhr/Jgz/cg
FT0nl73KpnIxXvAmkYULIQYxoRx4Vnwju+VAAgsg4z6XSI0b+23wd7Hg9oPvTM/I
IN0UcM72R57SZuZhtNB/U5gsLcDO3OIb0x6juZezYev6sy/FFBXxPJDdjKpQ5Zqx
x9hVpKDMeZ1esN9IXwPH4WF9ndsDND+rIckYvLAbSSAIsQzSFB7K/l3W++ewS1T7
k1UbJ9zqXT1dR6h8aXT1frMZ4PFwglfno4ZXIBw01eovMTIGTWPxcGVqMKn+O2/J
hypEDS81xIxEi/KvC2bbBrPPKtUI5+ujzvsdWxSR68uAt+NwR8G0WGTtqI65XJr0
aWQ+ShW99fKP1PXyuWG2gEG6a3zJJQHq7OPbD3bzQu2w2aBj1XsCmjWpqmogYg0l
W0RnfXeLvrko/ZodX/A/3IBtTK4YvOcLmbZHWMx1MvfKQpoi+pTAdNYASD2HjJBA
5cB/rP2eJHz6SLolfX8398wCJsWQe8Mt3Ha6eHh+uGjoYb1Brh9LrfYIvfZYtHME
cO0baVxg2IgsntmacjoPkbjG6ydDqqgcjM1Ek5nvtT9UhNKkDnscWHtYNqA+g2vr
BV+nbZXnloPCjr0NW4rSMWtP/oso8IbGW1bKy0rqHLVMsoNDrKdZE+z0JFcj6h1C
Zye+GxXeCR3Z8EOUTSWk5bJXAfrLeypetHgJWgBIGcTjwGCOnaGITKIfgSBKy7vC
adnabORZaTTiPFndDKaFUodeOZatM7ebRun7sKPqZLaJjQ+yst2tppa7P0ttkdC+
gONNNbNCRMOyFkyAs61sXXr0FhjF9qH5RXi/zh6t00CY7MfDFlLtyZaAVpFA2aPP
O4Dz3hFDwomGJcmq2gFJzFz3X9aeO3U6u+CqTcfABFv9tVW9LAOKUDcWoMhLFQ1n
OqqXALrJB1fQHKcwIJ9SQytLx/BPD9O0hBlq3asneeNn5gSwkfrtdbGT4P+SQlQz
N+mvB0fPlVVSYKRfBEpiOkxdwuYuHQ3s0n9MPPLI5NKAuKbofdnSYUlZvG5TpllP
Zst13lyrjI0zvuWb/XokZjpgiqca47PENwlMFAlF57GjpM5TziVezinB0iIrmB2r
fX8/FXb9HkR2slTU5pEyocy+TDBh3l7toTs1Ab7yqNIQ7AYTcSLRfIgmhSag49Ex
uJi/xNiqmXIxBELxWVbrtV/R8iF9XeJD2xzxm1q4hAJp8l5XbaJQO3QBZSFTG3aI
RuLxHbufQB+KQlqy71N6DP4+u+k3iG3R4wh+am6ZBgNkojBg8dXK1pyr8EFqORMW
R5OUSA5aoxH6EKnQMjKyZzqIqxYgNR1E3DtNKVtkNj++WmE2eO7MFHpvH2J0l2I4
+bQOcE/0sZ+PydKq80QyS8QYX1uudpYwtQaJEQam9091eHoegrEBcE2/Y4BkRF/V
H3Xn7pgb8DGXjQrKB4Fso/fflZa6jFIQvoWLqqcGXpmUkFJvxrVcfa9Kg4qZ8HGv
yREbMJha5cXBu2AEHhbQTAix/HuDYu3zEXDAadJkTVGTVl1VH6hkxYSrz/DWlVVP
N+jNObVWrPvXDCoCyvTItzURq5wnb7H++bs5Sp8l7iqADx9CMJUHoRJoAHrAjz+j
Hw2aCxDZdyZSwmUtcL8FRSEFe/e8Pi8lzrD3znp85eryGvgoTO0h1exiOpefgCoK
Ut3qcG7BqlApZSXWT2Rxk3Y0XsZVXlDSnfrlMsxja2WCYzgHEiDCNSheSGd5FmE3
QgewTp+U/M9/zpZuWivxFUaS/yNZv5FNvILX1rWomZKMsr8syHGRv03vhlqt55Fc
vthelucBYuj8/AeUNyDl15ITCbhgNMSD6L8vNpua2ej7/1H/hkCPCoJji2qtEvy+
cwqGMMpSkSy6Wg77ybmT318VwYQVo2bg39rBaJgejwJHjOzW2tuGg4k17adSled7
VHDCpc4lTgzRerI7tKQXDs5F0I3ArSGEQe3bkpBoDty/4i8m2gQbBrOBjN7GmQF2
ItT4be1h9eTOROk/hXb8LxXpkqBVpYgU/bGOHtnLr8w2k3TAl7WZMBa4b5AHszfD
jjfWS+e8uEmlBeZTD4kkG8IiQm3VZm+42EcKuOsA7MMf/0aIBzr1yJg55Qtm4Q8p
oyayCPcZZ4m2hdAe8w/LxGLK6IyhrZOVkEbHng0na3rCOp/kaE6M1ylPQKlr2nGf
B7bXQke6GBjtNCgdLVyA+NUjCz5tvNgIQ4n4FSUdlhP2lwE47b8VpJlb2JZjveHE
bCmEZKljZx8EPmM5KcR5piTrPQ6qqS2EYiqt7zVEAJiVqz9JhZ/3Sjv9eU29EEks
avq6Xwqg/Isd2Af41a3UGVdXwfhwaNG89Arh3V1vhOwGKUH+EGfeW6zhOU4x0rc3
RrM6fWg7ORXYLSngR3P3hm2g+epbrJZeWo/PQKRbe9iRK5vWDmbcCKH5UhyuUWvy
Cp9VZ5xMTnY2Qzoy6VvIGL13GlwUaL9C8ona3bmUJejgKAbp6mMmEk5yItmDQmFg
pvB2DcL0wMkVolnlhNTuEBMIqwECWkTTx+nQgCcURxgmjXZ7Nu0I5ljFlqLkvEAF
GGcaioo7RznDYHS54akz9U1MxRuOZSFdBdOdVNWu4MrcP8G0ZeWIiboZul/FBdys
/VXsO8TfkxA4KStnRryXftaQkBuSicecEXzoqaHzGHK7ZGuWp5FdSRoo+XqXZDsc
uSA2LZ3xUkbQPUipTGVZTg0VzQpKY9J5Okfj3WFwCSxo5puPYVh4XuUQehCYmE/A
N9ZF27F++Y4PqUYAt5U0m221WFfgT0a0LJdPIyfOdqx3kzunoIKaQv/55UR7e7bU
yRIVHSkmQPhoDm1vVLltGbTzrkVZS0UrfylOsjned+g1e9sjmQmf6FjMiGXf3CGD
4vQ133rLrxvnqGW2WLkuKSi9IZcn8rV3bCv4O6XrQCEDfK5w+dGMvKh6PQL9mZkc
xzVB+6DjxlAwVFRwc2Qf3q36lfl6ljEIkitCFhGjk3ROEudiuszjV9NKIBufaorH
CtplR8wtIlSdXr4aOdlpBnnDhob+4X4J+/pkY1ohcxd69kkbHnPbArV9elTq3mAv
X1/pwj4EioEBlXz8TveQCBX9o+fNNmfyCTjTcuQjkOaH3MfaowRv5zyiSp4UWxKp
JRXcOxkYazjYD1YL4C+zo0gqDF3ot8EUaA2nWvT/j9NrXQJT9TkVAtsQxd1Xn3TM
YoBwLHT8aDByvW53rpQGmV/AvAKLYvNvrYtC465AmQ2xRpOGjTfKT6767/6hXcD+
wZoDoAT8qq18LR5YU02mgh420134VSJ9ITFORyBLRg5liH9fzlw0YmU6bSwv3N+u
knAl3lZu9UNDq18VCt7Qtvb9/qajlPBNL2FRSM91yOVwzZXYWYiYVwy+2DAEVWyP
Ijq4/19pZvr6EghGmrR4sxuTTiPovHRHhiccwI2UwnpQ1FpTsjb8xTlM8ZK4Q97A
YgF9c6O6p2nlO+TImjhuGMGsLDSuJzS9CeCVHDsyoltRIDrjfcG4Vp1YdJ59HCJz
/gTW3C2qkq4PHqfz5X9/WBdYDdTskf0dHN2IML2yT+E250WaFqPVEOLxQFpRTOEc
iokTNe1yoNlLGmKh35E4S4pdBbi1EuwkVkErIzjPX+IESdFyHgszKgdDrrgoxu9V
P0O+3uK0NfyZ1jIrVIQiguT/S7rvExpXxjOSNbpfm4jEzmWvg42fBvZ6MyzqPzjK
Wz798VMsP2bFYZP5Ns6a86MLtIWyJIvyHnbzA4U6o0x+LlcpZExVRwYhxAdQ4OOk
kJ/1Z79B3aMvWbwInxAGD9LiQDOfdnRLCRYZEzrwiXx1p/sQtFCgp+QWORZ48+HX
hbg8sEaJPQv0zalxaHRvWdZ8Ml09DaFdMY2N2Nb418LZ1eLPzQfmyQ7a98vJQqEv
hDZ2V7Fk0aKgNXzodzK/UhbVuwrg06e2bISpd9K5/cUA5nwAkMGT0Tn2cuZQ3v8U
3ALvtC5BMU8PZb/3fvpkcH2ObDKPT8faksEIGaNRJ5MIG3oKtVgtkvKsVwBvt8ta
RbJyjy4vKdDnDDq/wVfkhY2koJ9hNdLRuBlU2UaaboCsY2400135j1Ma8ILMuc+v
GUttwShDFJLlDM/vW8MzHYZYcDp+PfuTSKX5wsJ8pWtC0J/GU8p9BQXRadxmBK/e
csEF67DMA09Lay2RvVT/E0tZgFRsw7d/Fs73ANGecNDmE5+xwCrr39Bv4rNWgOmy
M65wXkvrr/EhGvsItvu9Mr2OUjKD4cE24BiEnTOX/nH8cFT8KGe+iv2s6g1gqGJb
yuVHcYSdXOYQHDU0sMWjmC+nkGq9RwreujtuSoiTwO0e5M5pW1Y1JLZ8Lqxugh4G
wI6x/iabE3cXWOJX03J1w7AhCvan54vt0yNz2lLsWrGpvB5e15ObuiKVY8nkZ2Hp
0o6s8xGT2U5pXRtuVCMacnlWStPO8AxS/8NjDg2idohZIJnwmXdGi8vs7e3Z9P5o
H/qit6Z5sZeOLbLRIMq1hxRJZyOQN0I0JOkLj1pXDuvRPGcaSS8BV8RgYGDq5URn
ZfeOynvsaeatHRxYUUpBsKGlvrbbZqKfzmTp4YDSlxQrTYLsjnyeN/fhy9nAVXwY
/uy35CPaR/RbZkimBe7R9iCytvPsc5xTyPikpWrKCOgbLi6h0tASJ5fYzjNxpjux
PQSEeOz9V3q5L2P5shX2ZDx4ZcNgbWSV+qN2S+N+TlxOlheAFEGsRn0wbDvoRbQu
GxQ5blmC8QBDrJUhv1LjmfqkwEnEq+JE489DJ7jF/HRZJ5H8kR35AglY8xKnPoi/
DEyNuQndxFiVbsl1jsiEs/oZq0CQ7FCn16tr9dJv8eeo4V8HAV3tX3FPyF1pHuKT
5SqqlA0HD8wF7yLiLY4SnjM48EZrWKrH8eTGPom831SoY+c+N8qbmHN65/ZBD/3I
XZWIYf/Jc2cyJS/5E/trlzcxMNQ7HJJbCvN+mp+K7bSXHiR36SWnqFodcfmiM+kO
ulhzDS2sZzH579r0M1AxWFSYczyvanzAGMW9zJfJYwVlwAYDjZdx4n5vAIllwzQZ
kFQ62jqXt5a88TYOUtw41saOL7uImcq8gT5R7q8PlrcidixP3WiZRKoOcVNulIPn
dYrnHJfYNIFJR0fDfg/sZZOybrWfXWu24cCQBQ+MWRmcJ0bpoiUQYCWuy2e9l9MG
33Y4WO1RuXYD+/ZtdTQdDAvAV4Sdgm01KBEzFpyoTI3qw+1EAAXjIkMhdbq8/1WT
h002arkYkuzMvlFu8F/aqZ10yimtHEOXBlvmcGFSNq1ZC3aY1vvDXTqTce0wKNlT
/8wgl3bUraoat0uQIn7QXbtDjhXJoPfK/Hk0VTZNyfOCdyU4mgkPgiBej9P47I68
/+FLrvO/UMzCFYHPgsUrozoLdZM7EwPk8AlL/5XodoJJPUS8bq188h8za4GhHzWy
YFOxUWcVHE4AdPnWBnOtbpcQ60QlZxS4J6vlOkwDQujcB3aCgj70AK3s3Gmw/mBi
H64zp3EaUJCiRx709dVSS81W5Tysr7FVxNNtohO864YDLQyH5cU6eFAZGguZmwtz
NF3WDg0SrxvEgF0qUvnHCMpLypdHntof0XWIQelTVZDC859UKuIQv4n13gRHd91F
V18XaFJakuMX1/8HayL9IR3DyA//0ZgEjLiZ87H1nmdFwvC5LF26L/fAg+0ZF0kq
16Y97mb0V7TBl+kSvm/xr1DYKixmsKofqQmoFGxW1AFuYvop6KP+j7/mmmvCci6y
nGO0h0g5z1ahEIMv5wvwJbtVuPbPtOnto3MpcRqrgpBE2yotCfdmjvXHmMZDI7LQ
rD7Vb2+nAWMwEimRVnetzVQ3nzqKMDKwEzIvAZyXgVRpWb3TqHXhb779DtmFcw23
dFWvAUcCXHa9D96T4/bddsoLf7hce4+7L/GhJX/Sh+2Mf1Aw4Hu9aw+QemkeF5y3
m87mcHa1F8rj5LsWviJftCbt8dqynIUb2JKWHer2zLhYbwFKxuaDL7XamS3r8rz6
js5S3e9NO4wV1i3JLrVCB0G0aAkNvBeMTnQpwTuiEZDO0IATFsP4yUfZLuXebCQw
Hs9Rq2sFjwZwuRQyYhKu+7TKjiWlBlURaiitAXiaV3TppUBhTo7bDheTl8dJnfBV
36wy3TDXcTVfXJR894sLxV91h0uZhY4w8tHZuhWSJmY5d4iFRpPaPg9n5EzHk7d+
83FAOcx1+QYI+pveiDuV5Cbdx3xUGaaBti+709pF36mMJg8HI9fk5xlPUUxfB+fr
piEINWcgze9fdmStrS2fHhIA20xNr0Lwot2sbNtyLfDXV7Pw+leR+5TiQK0HIAXJ
quDYB9f42gSOyMr/GRZtGqkUepZMAsE+wBi0MDb+4T71qQqMuc2dfBYnzjekOENY
fLv6HmgkXb8wcILyipPGQuK4C4u/k13Xge4nHv7BPexvzD5/ScxC4HTWLEwPzvCr
2gQRQc6oNDqELZqtBFEk1csPVbcJe0sQgeN68+bf4qIMsjzgUDPlTbUka/2Moa32
sxxTtSubtgIyl+wS87fQ/znQVxW6JWyoJNZBtpHmA9j61zhMykV2In4T1kFNpKre
dKTep3O0jWDjSuE7Ujb+nDTRE39H0zCDHXOI90Fi9SafO7yt/VOPbAZtBeqQXYmp
3JEo5xX4+7ZMb/vr1g5Ti8+P6WFw2A1YwswWe3G002G0G2SVFEii7TzY4KAcXmTT
zh4IhcgxR3kVmGB4C757HR8wYoTp3qZcHjM2M9YMBfYLbfgwP5/IK/RhgpDq9zPH
ep1MhdF5jPHJeCVfVe24JI0smR3+IZZ+/59Woks4OIxne7Jgz2OPvwTJetxq4dnK
OBXC7LcUqBEedi3PdXwWzTlSEFKNdkbvLm+2juw/2p3cWso+c/ehs973pub7b0cW
oPqrdlqEsm07lry6yGEDnUOVgZ+rkz6N8ijxmWxDbsqvsFTKzCjQzYBZJf2JHg04
2Vv0ZXIPFReXxdgQrlTpEjsh2icsyo5plap2vaOhjZtYoYwcnnxCSV6ilxBO2lc4
Ov5qaOizFDiCFNQXV8MG0HMe0gSK22QIbFjAoXv2VRRApDJDy1auEtbuK6Q+kWL/
8QBv4FkZfJgLDrmxIIfRBfYuQo1TXM7V7kuw3pdJ2FXPs6GUhnzx+1wId1XG6Ghq
TfMfOdXJhXAWdX0aaGEwUsvmZKe374H9sdsP/MKK676z83sNU/tLK57R2Bu+Gsgb
wJJbwYy/1XEzlXzPQsMNp50/KFpfoxRff6CQ+lK28uMbfeAMsIU6VRfFcRVp70fL
KH1zJX9IISKxTGM6604mDy28rfcpKSnR5pKB5GMJvWGPPjxjx6yW/dVKufBI29OZ
lyVGYB2DK/s3OjFgfbGIXuNnjO1U1BLLFZ9+S8BdgXXstQrWXwjBR+XUBIN6h5hU
9dSPzxYH2WOhzW/nRy42CRc2Qfet/yXe3YPXOXhKXTKWJaqVG7BoTqMsKmqTlwME
sv/Zlk8xMf7nUFJ2cALXnOG15uvSOQi019mrKJhCvXmu8fgSkAiMnt/ijpanTh5p
RqvYT4sNjtctv1Xf0y2hfC6oW4tan/zKPw3fgRP9UooZYmqdosdrVBWfr+ug5mFq
DchxTiQwd8Lwx0baZ0mpIHH+dEmIuw3u4C/bud0uvZmnQUNR1b+cEXOnGGxIsNzK
hwXvxbMjIHXNUXDsxliK6dXFtci53skvQKRJMvLaRRd0nSBI2EJFElyIce9+Blup
HY6rhBCZOhNMi3gUDpaPwQlWMLtj9gAaDD3UJkBSG2PeiH7WLo3bEZaqEwFEGL92
dDcvaTIzy3Nbur3qY+AD1CWtaDurhBWCzX+yU0tFoQq8Anh5mEMjjP6mq/Yzb6Yo
PrbLM6d9TeRghhId5jacB4bkTB3btxmOu89MdZJDs3zEnzGnoEWET6PibSjMhN8r
XKH7B2yB26N1xCYijP9jKH91FAtNaHcM7jdWqow7lYfUP9c/msw/e3zapbQO++15
7AHoN51Tl4WR4+/ryeHfoeBsRJKmJT3mWWD0vuMjoBmSE/bmrSMPdz8dIDXmHTrH
RDqXBSyRXi58SHFVQRNOUTqE/3yo433F2hNtSvzKggY1o0I/21UMw8g7YvymSRvZ
5H3wOMSPUukqmsDWwC1dYHesCC+ee+LghAG1dDy5WohBsNLpExf5v1T2d9YYV8zA
otHnh7VCHrDQHepBggSQZBpn5T2qKRZxswup1zobEcCBjLkaPRcBK8p/yUOP1aVQ
9B0bgh4UU7PUFpVby6SA7d+4eLYPnGVrRBAQSEijneMl7l89XJujU9xiX4ULnx2U
GuLSU/w4h3ub48tEJ+E+6bWWthjeekeBt2TwRSV6gooSlmrM8DnE0o5s/RsTcNYb
eBJZ0yltlLDsdhpcKqpkTH1dIuEXd/hUNZwdbOh4vxxyrJoAcqyTFqw8ckCxiHeQ
1/TeneOPgMm3iGxtJbGzUd3ZTeo2Mmji8E8zVD0rqTeq+TV5mgoD8K0EYksUmDJy
MYLsL+rDFdn5602+cLdFhj/BbVfwtGMo+5BaN2keeGVMMlqdo5yA/XCSBDQb9Gcs
YS3bzuf64nBs81WpCY+JwJVAF0QURJvKvkF/Y2Z0pv0ntuOCcjuQAlYY5N8IY0Ab
KyLcUnDxhvPRP473hau1Tl5gHD9DZ7cOLThY0qUJbXRTcJzoJzzpUTHg57aH/KvO
yR7TS3YvYL2hUc/m78R66GaCUm/J9dKuuplC3VjVV6Ea9/V3LeyAmp0WH3iCRjxY
xLyEgJpOFiSnK0D5jm7vx6lUU1etWMltm9YDIZ1weK7pfnn4p/un+LeEJtpe6L3E
xmRKfI3xSj3uAGf5ibD9gyWy0vYj9H0iLktOflTsSt5NCPO4ZIAaM83YFHIpZNbW
iaQCOgKMZVkT0zmuUCWxZUD1VMXbAbjElnXEFxpLelZZl3r/remOs66YrbuA0gle
gC7ZZ6dBKvJCLhT+pDSv31oGKBWQDFm7IlQwmb0Yi2RP4n4WvSFJTZGz3NoEiG7m
FHJ+mDK7f/ZSmHBU5DPQm8MBIcoGinOewBF+4TVxZN7ml6S4CkEDfi8GHlLye5Oc
EVz4lVUEH7V+Lg9bBFBxvpO408Zp6Bppc7wtkNMboIf8x7Il86I8B6TLCYsKiJbg
dTprocTGSZzNANxnLlcJTB1wrCX10y3fHFEypIUkYCRnu3f4z4FjGdQjzfw1U4v2
3HhycVCpfpcw7Ko006VqrU87r3oUhMji5yPHyx7L4qEQ8jY8VfWQDrbxlt5Myjzb
V177XgSjO1XDH8lZK1DNRNuUoyhQS3msPbESpwEKk4WrG+XKb+di+ZuTyiDUZ8PU
wcxQmXfEJYhmzb20PmQAWfM7Tdh/r+g/im1lVLpm0ijns0kte6kPf8lfuG80B55g
2aHLIOhkHfrWiZck77vS4Bh1S14MxzU3EcMSaGsPg2fiATsTRbIrBlLcrsHMG72u
VFmfh5tbGpHVGTDbM7tKtw/XJTlq+D6gRFidbUuiuB3oO3AVpcnZKLNKfa6bYp8H
KfIDOL5SPpDj6r1ZZh6qs2GGuxVEqeN4K/OfOYFCxImCE1jv5aV2FHHqsuXG1DUs
6plW/XJ+L8E4gcy1L4/Qr4MZLbOYkZG2zE4UQofttVUSvFmKOJRklPyBVSiYuvPN
Yy+447XJ8gQBIZtKK0eN1VWsHVppF0ej0pmcF/z+F6f4nIZINJ38iBU+R/CFeqzo
Uht9i7DD4vHoYZpYIk1SrosjkGnUtvuA5LTEVRv2b9nh81fMWnmcn+/KryZ8ney5
hDPv7+8NWyY+p+olvXC1bS4CeNs9/v/W+yuPs6FedQFpIKAUMtEjF6+xQpbA2v2C
OHHMz3dDwWPSkv5gQeopJ6ex2pHNyWljmznlP/ONZprNuGuaWoveslLdxTZtZG9H
EgOh4SnpYg+ZTF9DjFgnuYdNS3Q5GDDMCF2tMB/ygzKUj3+GEDJFgr7K0CW9OEhv
zWUCZ1PE+pc2LdaOBGyc3IzWGOnBUiwhaPXQ6gNR9vf5Fex/Pt/su/0FvwAZ+Z0f
Sz3VnCCdDM6NJDWaOIEd79EndIaDmdtAbd/tqSYXMKOHC638Y6Wbpt5pYjOF+RfA
/aqGs46sZ9DhBHu9vsbXsJrfvzt8IisLjy6yKxw144eUEakV/jn/W5zFaaA5ilYa
0CEqy2UYA7L3rxw1mvF20Gz/tfMMeXa4HjkIdQr14svXAXvQnxIGCCnL78BgWVfk
eoFbi6wPYWgSU7ftdBn8m/1tltr2JXntj+lsM+g7wKQTEN8mKJ7f+7xI4c0lMT2D
3F4TL7cLSMGepOtHt25kMe9M6q7IpEBC0dYFtX4odgVe8XW5Cj9cDiQLH82dOZFC
r9hmL2LfdAP9UleH2dj7HHfQrusVXLF/33fCWj4dzg5+RazotSNZIMmfOcm4Z7F4
ZomRo/T/Dd4Cjt17RWSBym9EcN6s+azQcUw+AB+w1ojbtXN7wYDf+pzBworx0j6F
87qfW2L3/e1MrWGSvNnZWO2aGsu60zY2XKl1E+OuvvfSkgZ2OSz62+DbxuxtmVr8
nV+wkpm15L02d9xM0S2IRUCPxXvKJ+oAsjF75aicEw6xqQNSPF9uBqF+SPLMq1OD
RA+E8zLir5lu0vywtzpt+TVNRBkvacNebukAxvdOnSBvWKzz/fT4+yFZBBUGbgnm
gXBEdAJiQ11NaxLCgky5Mo0xPN0Iem5U2rRdgnZmsPatmbHPCHWu7d2IO6LDGlIZ
Bw61jJ6VuQGJ4RNKbN4rZzOYC0h4u4hatZZPnQeuCfiURfgpSpW5HK/PXvL4A8xW
epFgMGQ6dUO1y3Uc71PmwvDU9wBJTPcp8SGwg9OzlavS7knTrux3u37G2T0gBXoz
UqXmAM598YmfBbzFSGy+9mukMIHz7uecmunUnxuSs/5lGsCcq9L2ug5a8/nQQewJ
95jsjBRIED3gHuN+QryX/i353uNcS8nG04TRThN97ZsPMazIurnksUw9cUXN31nG
AD2qaHD/4acbZq4sppLMxBHsHLMm0uplgpNk6ww3BQxggOeNECgQdKoGEi44qi2W
0YO2WHvq9IoQa+PQh2Iu69BLLAQFl7xF6D7vb6eVbuwBbw0URQJQII+vbDG+9eeC
GVGYIVYlDTtlQHG0q4CzDybmX+3cV8DQUPGhfDQnXs0hIAceCRffwVhY3qFoGfa/
lHaMR5rgDxygWyGj1/+8PU1u3tPi92zYwUZIX7Dbz5+XUXaM41TPE5N6muFbM1PT
S9ge7mfOUCVopYtvkkgTex2MGAy0OqP4HVUHk6kUnpP86a1hREOqAOPq9kzFOHFe
P8fpcNd88SyIv9ParQyx3WPJFld7GcIBpllg6ktIGmErmzYZZ2gGHo9m5gavWAu9
rgmaSVQhyaJmDTQDrJ8okurqh+1CyqOSWHYaGGLeXztb57ABIfoKLPjp47zKJ0q0
mhvlLnbCVLY1K2MTi/2O9ArPMJ8jm7SX60pWvA/YcGN6yCpJW4+Y/i4MR57mHExi
jyY5XNybHFLxZSLcpRHwy4r9FI4meGXz0izGgoMWG30JRH6Gz6J500ShsMLz5nF2
BijZQ+fevu7wWAl2inb/5Bp7vZZARgYTHHpfO/KJpFozFusx4xfw5Nm/TPeHwKSy
/dm9l1PgGGQQjwIBE6PaJ2jW+dFvzF+ZVZFVTO8a6VFroJd6Lp1pmOr2ahhrPYbT
5C1J73zip5qzFPbqz00EgI9GEcH408gv6qXvSrHZWP7765jYA66L1LGlhqU6FZxp
xXfsC5KaUfoDgaC6Uf/N5FGTSZAjliHF/T87TfWvkTWjQTcbuuq72CHwlHYJS6sZ
AfpSyhZnZ42olHXiMnL7gjPg26XqscvAZ9Tj3jCwMV+JSc68zKb7FNRWZ8HdrVNG
SQ52oky8W6pJVKyCLYyoBhO9psccFXvRTlXHb+EQag2d+gOkVkSuMD+VHGQBnzj4
clSaVRHMtM6YqFpFjKztrFK3xQeOi95TOMsW5cg07JEOall2EGpMm0UQi1Yb6m8A
rmAh/cTAjXVg1EjrxemfP7TlJ34Gx+JgELYGZGKR/8cImolAA3s6J18xLTGZZrQd
SEWsx1Zah7EeD+hsGPyyaNrVvAbyjBGLVg6oyKiz0svHOhrsz5VLVLiKjQganFUb
2vMwfT7mhjAr9/F3Y/nWWU8c69+WlmT4M48P0o8BGsk3sAC/AwFbBhsTevXP/xtT
a7uDBlLqxjOTWdjIgqvWVflRJ+aKyt3vpmvUhhtYo/x/msOe98DWPgg+Iyf3+Qih
Y5OlvdBXqI5U55BpcOfdo14tw/5aFhGBeIt8+d7sOGwW8oPvtpiN2P4G7ZN52RC3
BwLvp9Fpg3M3zsXkPz7NrGXfQcP2Lh1k4PTem0fNBlA7lO/OaUcycsL7AXTn7/Fy
HZnzvAJFNZmx/vOXcoO7eHsgVhYH1/yaYnsfyR7vzmj/FzZbV6fgmoAYhbEeRMkG
nqTQiky00OS6ERDZNCCqu4P8BE0IWv7ELlKTJyAdmH5aAFBE+cVZJvEFC0VN4ZWA
7ypNOUDHOYAG+kVKD25bZAsvYsEAHMJ/UaNcQ0WvA7eXMGhHwv3MgZJ5uZB6Aa/t
7oZ1TwKMbPl95aILX/sI5lUqs0PnSi8xNf7ZzVHmx5RbbVSQKWPGUQINZk+oHmLR
MVGHcHHasHmXKx8ITp8fbG4NktcYtcAPi0WKEfHotGM4HGjJy6S40LlLdPYMl4/I
EVy1wa77A66kkK+1ZRJxamNFypC/yrwVqgjs61fihEgkaY787861gulEuCzdT884
WLRZ3ECZIjlPfH2g0DSLHNK86K8Micg/2B/UQtTUFXyQp08jGDBqLcMWHc/XHXSi
kikmiL86ozly93/ds7ZzPxXAvZjJact0Ssj5Zjc/fptIU7I86u9KYunjUlEYqzPx
lMhSfrieAawYcLEfzqOCDpgl9sIXNdWA3n3qm4oGALqpQTZoXTt4aKmVrIUeky1/
ZgPr9I9eJkugAHb25nc3PM4cXd9kIShi7ilTuUp4E3RTbYWcbITpLkUyVJ5nM3/N
HknPFizr8vRcwRnWE7H5glY/tpurTWq4rci/NFC15s/gEe/4cW8Bhd2RpRQ86AK/
0j7ewZfEm3/U2D5Cal2qBMBa1/nWC5MMSnVUhjl3ZLkV5SQgo7M+BeNZ0dEsoUNl
NINYpJhUgQPqWp59jE0vJoAzb+/qDS6nJHOt57s+8bqBqAsgfwFI4DmOjWXlEcan
6RCBX2PH4IwpAKwLiz3syIum5wDb9dvoLtjE4qKEQPx7ct4RsXjRoNlIXE1nIaVQ
EmEQLuuaAJtpma/BvB36GjCutodTLSvqDMxgPM2IDX3dkzpVHBelCFkHmKQIazeA
Wu+J8YxPmZUDF6NnG/uDcm73i7R66JbJT59FiUERKPdpIGoViy4tMzQuJKx5ClTl
ZCJ4E8YypXVXoLEpVb3Orkzr+eu2p2RPU6Kmn+KO5VEqEecChIqy5Y9YnBPlvjV0
LzWvehxA/UHh1nOOiEjqtuo4X40SGOJcIZXk5SoPYGi67hE1E7BaDP8jaPPG4i9+
SH6EVsfrA9xY0uy4y2Qy+D30A4KtECIYOHp5mDI/VYqJbM3VisrwE58oOdNZkOwO
Gb3GJbnDdGYU9RB7jSG3rX1KJulRpkM0X8tJXqANQt8ie+aUSOpudFl1PUwk9uEC
msLC3NjWhYpz2pdMMLxy1RJ3QdlxJJN9Sn03Ww6PC5FXYjLXQcGWDFAZfpHcrP53
nrT4pIsb2DtnHIF5Mkri8AE7ftGVA1h+xNP5VDHJ8JjCbmBa6gCRabivghaSdrjY
PXCzVsh+mKJlnrJ0gM+AMFom46xBKSpySzk5UrClxFKRwNL6ANzb0KJnPodsXNZK
Vjfl0hzpXvtAKG17kO2MDahbgv/BvW4icT78ht1lLXBjZ8jTjqBWE+L1cySPiRlb
nKKF1L9AcTeHdyKU3mPV1rROkBysCRydmfxt7qiyk2skPgGgi4BejoQ8R5fewONr
EDYWYmsZ6zc8ZjV1B6vMKvlgxP5x9svqDHfCCJf40YzB9emcTVz5rGaTmZjwX3nH
0WQggTa+pSjG/gZG59lhfCgsWcxiaMmwpm6+shSMWy/M+5+r+sVhjLilL8eCcep9
InvJHf88+w4pyKhPwQjtgBAIvvNhh43OaJsEt3FvZyMY/LYyvEmto8rVy+RBsbEI
RRRNFzsPLHz3LYhmST+CP33qmNtGkuUq/I6YIf7Yg0xJe8eyukUCdWtUBmjlt56u
K0eMUk6F7MxHstcWFvPR0H8uAyaJwTZQZPOyRtCB9rWKZr4CE8zED4jKoqBm+MFZ
rC35Km6aS9NrqqB7CZj9JYlRqfywdY68xMPTWDCy7p2gEC/oOLLuCbPcKcBIhGcT
vuZRaIS3Fi4j8siBrVhRZQ5YFDtIM3VC4VVBag5F3WH70XL8Wxm2Y6DWvaBiGO58
R/JzFVNoYOduHR2xJGJ2MkzlISaCXGwcX/F1tiqEgKkPILRoNYsfrv0q7mbPH9cg
mPbm8xs7CEXxo7TbdKYY4QDDCXlITgcHX7sHlPqqcAIeWejG6eDsLRRycXDnGTa6
XYnKsdyOu2MpSV5aQcI2HaKtz8Madhp4IwxjWgfesGdACwOxHnvWV6JnhihbiiSQ
0M3QexcQyBRV9RregXAs8I4Z5k6hXvSXhKiJhUK/qkznlLs4I/f+nop2CrqtTC7w
Sv7S5V9zI/gJBhAVYqOUsB4/ZUqjxxDaNpomhVm1/p1OkgAD85ksyK+l5a8GtGBa
/B1WVzi1bWVGQyUaR4mZIZIj3Ng2jj8JIxRr2r+7z+JPIngO44NkSG667Swiw+Ss
y7vO2qDhkVCKfLnZUgn6GSLMah1Zo+/F5XAKOknVAjTflgbakI/SIZS5bWEEPPxF
XDdmRK3NuEONoStf2xhu0FITdKUdP8+ZgsVK47ax0SCI8ckGGtBCQiJOoyVBdlch
UuzEPgdPpvMgBIyocx2/LsrImhh31F3xQGz+BKrtSe6pHx8wsFZ/oVQBdpPhjKFm
ePv5SoEJvNCzFA/ZHr9ScPdhQhh6ZYWJbelFBzbPzg1x27srhSLkLgOOBwjK8HBx
3g97gLvBN5y3TUHXjyVZl9MFbapMrMKMH8jfCrgx7S1UODigyFuecTgRj98aWbbD
42P6/yIHhXuX3UAZgYRqycj0Aj0wwZT6LSjK15OaTl8V7iI3poJf9tivkefl85K1
ESbHR9j+LdAeYBUTdD1aSmDQDaA914zBfyyaLmjCgNwvrumFi546hRtb3S9In/BV
8ZdQYF+njeUWPmM18wcCK7eKO6Vw05VFZ9EH/wMMLUElvl1WcAyb9R8ocHBy5A+N
7rJK6yXi+Adyhq7mp7HX0lYSkjZIN+vb6ABesWaiwdRnE+WK3oa8qSmF2fHImiMP
KvOnjk1b5F/+HD0PpspUYm46boPUPF4xVFn9sAQL/Rs2p1tkR2ULpVm14t7BIF2h
wKPrtYGjhd+u81/V108oY/PBrDOQR3bvdkUNX0GrSGXce5KRDDTa0Uo3eiw1OCyy
R1k58XJirw7ObANYAz0XwbYOGCPee9ilYlzOfSLChmd220UYHZMBcUkLf4vdc5ys
ujTvqvuyqhdS/gj9vOdhprYm6Cj/MMQZcMYgg1sDx8p9b9Z7BTOa+x7cV/A+kovl
2KnTjJoUuWdhGXTY5pZWbPL7AVG0Rp6pIM9QT3kEtDOmUBHm/qdlw1HxNBOta1Ll
M0/H0fGpmX0Ptl0j5VNGZBNNPoqMrnxCtfE0A5F4tHvavRoIvpDPG4wp7S5VaW4O
lEqIwxxr1q5KH/QsjqfI91xAVXbJQ8rGsZ0oN5GgAwza4I7NGDGsr/6cqu0mK1Q2
kA4W46woZge0r7LJV/q3kbtpJ3RnSSFj43NvkEFrOhC81Lib3/5FVi798gDhfH0n
0kjtf2TqN3Qv77NUnsa9Xh/IO7unoeP+zTG7EjnfX86ZnvGWNcpntMJc+0PXU1PU
zRfPYDT74CoXfc0X+RXUmTBCIVxb5eZuAFFDlR0FC17Lz0KFsS1JWJIytfx6GryR
nCYHxP1tvB7odBssakgjauBDP4/KKRJb8/J/JV9MHPPBga0QYLo33NyjlG7vi2TD
8gHMFl8p5HCNVy5ldtDk6a6QngUfIPxwfz5cKY0SRNa/hbpD0GGVmozekVafWtGm
az0cjae1rxYhygwrlw7i6QMy8fPZw66n1IzvpWz0A4xeik2lFKr0vvmkYJ15aIkS
omoONulxFsQz+CiBGBfK62DLQ5VZ3/Y3kTfXBShPS352lRj3GWhG4ywWpFDLc0uM
gkY3MycdtCN7x75573FV+hUYnIPvorRbdqX/YANDiqMRFsj/KyUO5mQLppNApRd7
jOLmGv6mPiLgdX28pU3byZYpPeITQEmMCkagJo69oa2TyoacCZZLduVO09welu76
VHuRlQRGF2bqfyBBWcqceaiUtCdNzaiL/fgLYN3lZrOhOJlCuFsO8BmoXEME4pHK
h9iM+IbfC5VX4F4gvcclQc4uIICCz0qFlDZ5mwhHE8Ls/UCJfK5SB4+xy9j0+JXF
ee9GFo8/KKb8TJvbKQt4z6ojqU62SQmmXx1gQZjYv5QQDFHTtZT4M3/LwtgS8X0B
P1tlQ0b11UxgTE7u6RyG5GmnJL1FlYmuYyZjmo7oN/uSoAcMjeh6ucWam/aHNFYP
FdURdriBcq2Hd2xTHY6FsePjpYBoEvmZYjAtAt0IBOSo/YIrsarBXA7T4EfLcuu9
sONA3WVRa8l25eHPfPVLMpJrGuBfebPTG4x5xsX3X6dWE9Xf195X7EboLgIZQhRa
jC5M/vfBC+G2O01gp5z7UacEwbcNqjX6emVfwuXNt+FVSDXfUz3QgkC7EYAa7gXl
AAR6WTPbg3MQdkUg8eSdGx2xoqHGau4i4bLeZ5OnrcNerU/gyJr5TxFwt6ZHljon
wpZEErjf+IZ4Tq1kGESBbxundmkTnPrfAvX9ByS7hlQv/2MBPOl03vRTUPiJOyz6
/BX1ifXHyUmbQDEz/qJ/OrQJrqLTpv29umjDCbeoYyyu6LBk2Dw9uYD8kObKbiWq
mKCyVB5SLNekw4Ci2aV1WYtSwMUH/CaI/bePmZOJycx6FVKuO05cUCr/gBBDT1Uw
QFD18+he+zNEUSFOMM/mvV8W40djwq7nmrIXW11kjfRN6j4XyL3R+H/9JB/UMlS4
YkNH617CoF3g/hxUXFOjGYyB/pGQqbXZKH0mp41PhGSCGjJ75vSZVyMnHyZptwrN
a5O7qaKY2nBrMvb8TpXf0SLAK/cXTUelTs6VFZEKOv04WKClF/1IYMtKQAaaesJw
ePckebrrx6780CYbPqzkyjXBNh+vvAq+34GI2ch2pX/ooPx8pBLLaeIi/bYXkSfr
YARuX1cRbDpqYkJfZuoIAFTp3YwSNfXNmG17YN/u++iEfCBE06/l8t6P4BBp/GvH
8Hdp5REiaKRDKmP8t22vBGlwE0wxs89mc1ZnI8ByKsimrfh6RJppyOcfH7CdsoTZ
EJEzdEgaK6gKApovaIwnvyeB1gxMW8OKhm36MSASPOEgtdpsxacnfGJYkZCiTgIn
fasarDib2M8Ia8eo1BoFoOxh271dwwd8XZXyqnrG2J87W++GsCsQg4pze63CErZS
RLkfVzvviLsfwcZBS4K41t8vDaMpFxtJOGINSL+i2/achuONeF0EgyawFNyooDLH
bbV7YyPEFgCLahhf78Qr873jyUqvz6UFmu78TuPG5A+u/1i6pqFKRaJgbrw49g+5
tUsYn2Mbt4nP3xl9P8vOV8K2aigXnVrenk/hEumITZKzWRtR8iAraJKdHECVrwXv
umR5KSpEGfyJpnnADIVFqZ5n5srzSGxWQ9y2tFN815J1R8jrPHFQyrxVfypusSij
ObySr+V3hRW5JGfQIUeHaPGRhYasoR4zgN+uIjTKOnnq9GZX7O0k1dOFa8laQQZR
TNGu4u6Zg730QmD7nKSY51ZepUYsDAv69TmdqjHklG7irOAOvQNgopUi8/dcLIMO
HI5byc+2vQuZMZGMi0IdhrFeq8wKew0y4+RrB7TKbvbWddefO+cRd9ynodP0rx1D
j9FSBLqAPb+81WXCbLKSw7ORAwNZwTI3bPUfFziYwIgQygzxZm07VhCUCtXc5R+X
6FNsSSeYbKIXOyCDeJKIDFUj0DGt18m45aPfjwUQByvUS6PBp7n55YNtFEqdOwLR
BeZtWPpjfSmhr9u7Z7aPgc35ocikElrV+Hc0F1VZoqS4hdNbp9WF/nRTP9ZWCZwD
HJ6wIJ2yMTvai+wHHKeymS5JtKJRBTPYpdpJWNII1uQNASAVbQnChASRb+62ASP7
EMe+Dvbws92KGd83xzAuvvBFN/VSF6YG40UerM+XiV98xJotMsY62h0bC4tr3sVF
sdSNmMxTuIlv4pG+RCLE6mi9lA0rO3R93ypCwdiJlBRenq9wUSe63Aax5KXVrtVb
OlMb9HRm5Jwsvgw9AOIUpR3UmPt+gZ5YQ+VP4VwFOdr/UXq9My1Mpk8oie+PLpaM
Et8dLAPwN7V5c104TLNXu2UhumCj352AicbMceFlNSB7qF2iqx1VKO66o6gSzjII
zOvMrJeDROg8bblK5xLTXJe5/3aePFKSyyjg9l7eOiATIyeV+4S1XkjNmwcVP0Oo
SwEYpz73NuysIAXUS/2UkI8oyTyvo449gdOIzYEhnGk091blnGf0F9vTfXAtR/Je
KLKDxIu3wX+vNAQW4a+N7UYm4QakdWDcgnCJ0+GNVe6FGV368Vm9RNB6zAYz1N9h
YDBIXyof4ADJZrnY1ckStu4646unq5sxQfr4eTYCrLTkvnspQbxCkqnQR4jTSG8h
dbpcvUfTHyx2o6RbOLR4ukbOEN5L6kANH8h0oKihiyayQv/PvrMXoyQEUuqc4WNw
qX5YOFHFcyr53WYbtcB4X+FIbuzxWTOGAVa8ljlaTybUvfyPCo5NPX2oTAUIe9O1
Tqmzb+Py+bKssPkVP1hFa8RV9tzAL5DHiOm2XHfR0VYasSXb0LoE2E394LUhWZaU
nWjFfNiyKoCZrkUn64Lg/2GxAC9IyHESx9wDV/V6L9R6vkkFwQyZnrPf0Fdk1zU8
Ffhpzsi4EqO+5DEIHFRDxvehuh7qr3D2SDuHTdrrJkMMurYjvS+mlYdzAIFfOTJl
fhQX5ip8KC34yy8hfcnjiQX9arSRdUOljwbfm+xK3vU+cmUDwUiq9Ny7iv5k0zOO
7ywx+9eJDkpZRihLsAt2egh4OXfAuz6QcNbJwmmfffmxRUghNQt2rJwx/iVi4hT5
blUPOuufkcWuUKk0E42iBAfuDOiYhyLYVDHOP+oEmsI8lgFrPHpKwWcT88k0MXK4
p6/LTa/IlTbFYHSEbKI77qsJAvHGl0tWpujqob+lS1yzbkZLgxgIz78Cw61kHXgy
qfLO0+G1SNORHH3JXRkGl69GFy0FotJxOc26kSz5Y5NDcpceVbtxJFcOnrV3FS3q
iNFH3GcZO5O8yLe3cHel322scxhhFBtPr2ChUBb5YZmdjH/NS8FmQuNIKGvOp1Yn
SKEqh+yomCObKQkbVoLIN5BRJa2kx6itbkPyvzfsP/VINMx9g6ZJeqZ2chG0Asqw
iCB+pdKoo659s7Fux2HZBRg34tjyxBNnJ4bLYzOlUSfVJIckuN4Su8MPX/ajIEEl
aYWtHgLzDtk4Rcy8ozSel5+gJxycSH0oha8Fd6Wz+Y2AGALrkO4Zco0+tXRNkq0w
GwNQyAAW6k8N1FLSpjfB7nzjDWGnF6MSFAOLb9AkS8nq9UVUsXecootuMelnl9tG
8JhUHHYh0rwLy2f06gF9hH5ofpoyGJVKYb3mwyii+gCkAr/eAdiwg1VrAQnoaZyL
cvB0ySF1I98jeUUWlg1b06gXiNbn5/ikx2atGy5yddfMgFf2AllC6uNtDEz0gQU/
O7O4xPh9oTIFn4yrglZ3efOtSzXa5sQtNkT/Yuu7Pt51vuAZfMonHRZE1rU13/Wx
2sGzXWc5AivA3/v7UEjib9DxC6h9YIeEjYQpeSjGA7TWRxg5referbTfWqaFR9KT
WxEE4nHZnyQxf1Wwd519i02kRmf3fJBxokijlEn6xU6DhIV0hVAt9zE61+ukM7ii
lSkW+6pml7B848Zvd5Zn6ZwOJAPIlA+Jy73L1E/fniVvl0vnnkwjyTmL0MGcT57l
urLKRfe963xElvxxQSYtfyQtqBp6aMP5PWUIrfS6epNSSpsKk0I0oZpvTxANAQTc
3r+0FlfBLoCP1x2cSkPjjxOdenGZ2lk1lLD7KVS7cVB8BQcNEKaHPlyj8EMrcEr2
6nEVmNCpLxNrKYgGOkta3RMDjCY5RVzt7zr+SVHyM2vKwgcNL9P91yKFEqIKufBM
GvZ30tqm4UuZmzUEUiypFUGp79oss6deq4g3Dp/yF5/IIlV+++HssegKuZ49JYRA
HKbkkVF0peBwnggYO9tyrseLwQrjdAp0kXxlMq2bFFkhuBwlQY7X1WfpMdyO9dVT
TFtRxY7FvA0vox1YiSCejzVtOHP30bCZZmUHthEwSk362Co4uM4utEKtRk2ghjJo
/YYvNrKgUtDR3FRvXI0N3Bx5UFgcnEswmIsPYXLJhuVeZPIMsKccj2Bo/KN4W01i
vZCZFli56g2FYqQFWSIEvnxSDsrB/7Z05IXQMCQCaVQUtfpsOVJz9+0VjidoHFfY
gFZzBeTWDtI0Qosz/t553fTJvw4ubsAU5mGec9ognZ3rswM+vGJhFgMKgfRKCZdp
TXs8c9lxuLr2mQ2Gr67okDyoIatWGkIOG+blPd/9cDkkdS2DNpJH/2+8elyeW6rN
1BYzxXQP5vWhNK3XYycgptWVjgSfuu6NXieorqpuKYGnUCbXi2qFeGy6FnlN27sz
wWm0x7u9rohKpucEqfzqncRwAK2WsJBCXTo3b3K+EPlYI0wt8zOvd3H5RrBu7K/m
//pragma protect end_data_block
//pragma protect digest_block
9sxJ4X5ws4ARPTc+kiQXoGLKUfs=
//pragma protect end_digest_block
//pragma protect end_protected
